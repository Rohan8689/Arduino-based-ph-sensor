PK   �}XG��   �Y     cirkitFile.json�[_o�8�*�����䐔��m{{����
����$�V�����[�)9�m�.�a������g��sЩ{�,�Ӌ{ݭ��	.��[�j�J�`Y5��]|���6��l�G������n�6���d�(R�I�G8���(�@Ӥ�zA�������'8q��F|N8+c�H�"��8�E��:�2A�Rq��<6+��X�$5�y�d�E\p)IT�:���iɘ�EX-0V�Հ�:�mU��G|�n�Yw�<_��<�0hC!�2��55GzM 呧�"��Hy$��z��%d^db$� �?@���$� �?��;�?�,=����33��|,Ѹ�)����k���ڱ�@L-13��v�#q�~��~�n;��'�~�c�K�-�E�[-e��1�"J�"��^V�x�"��T�BK�u����t�/%$N0j����1j��E	?j�@���0�~��A1�A1x��~�0������������������Q�z}8�w]��k ײ�tZp��Og�b�t�v-�O�ŵ���sA��U��m��}�jdA��^�0/Z�-�؋�ċ�EK�u�����|��R? �~L�@���0�b�����)�A1�A1�A1�A1�A1�A1�A1�A1�b�E;�x-~l��r.hOjq.h�Z����I�)h�������\�a�Puz�X�*���ԻmW�.��B��1y�����?25��ƽ�g^p3;Vޘ聙�#���13�o���f���77OQ��w�	3�)�"Ε��ǅ�;;�d�9i��B�ޏ�k80��=��x c"� dh���oB����#R��l�UW��f���~o�2ضF�U�m�.�-Q�< �R�޼���W�ꎤ$�(fu	R^N�s�t;�CQ`C�ס�y��o��T&��P�V�ڡ�R��)`q
谊�����E"`�X$��E"`�ȰHd'��ܣtˈ��J�|�ܵt���K�h���tK��M7�9w6';��j��V�F�ʖ�.x�����^��Y��%�z>6�����pЁ�r����O-3��ԲS�O� �`%`�m%�J�� +V�X	��J��4 Lͷe��3����y��������5��H�=.��O��z��p���B=��ܸn�4t���Gݧ�ToS�L��\MT����ҧ���t6C0b�!6�!nc���E�iUd���/��lu���c|d��?U���@��ڥ��J��n�����̜����ƞF���v4�U���~���6���L�O����m���.JU��\��}���Zoi��c]u�.�n�͢�T�.Uޯ;ݝ2`�mǒ�����Y�����H�'bg_)�%��x���H��Pd�%B�(�$��,�3�D$����z�����00ٮWM>*r�ya�v�ѢF���ꮺ�֛]���X2In«���3��t�G�:M����<��?�a����yɱ8�D�Xrd@���%�-a~ ��\�=�����xr�(��#{��35�WA`����#�}���C�d�f�S7�f�3��Sߏ���G���#}���>���ѩ�'Y˶.t~�N�upq�~�}~{��AUmN[)U�T��Ss�H���JBA����?.�ք��w��Q���EƍDYD\Ae����4��<��A�ο#g�$���%��&)D*ύK���9Is��{�,���p���I�0釦e�T�Ey������\�i����_�O��"��J^�Vu���P���	k��$��FY!d���M�s�k�um�v��-JK�2�"�	cɒHj"#�MT"@g0��uݮ��5��(IӨL�M�`�!IF��*x)6����R5��r6�ڦm�����5�e#�B�w��w{B���e��?E�W���cHC",�Zπ�ڨ� ��J�8�Q�-HR�s)KYD Ne)���� ��8K�%f�YN#Fs��DIA�9�I-�"Ny����r�`Dꈨ�@���GV��D�?Jb707���&U�b�<a�4����up�V��J�����q����9;��33�٧vݍ#g���Vw:<�۳nݜ�&�]n��q�oPT��;U53j:�Ԫ�E�iW�h�;]� 3X��0��l�vy4y��Iz��R~3$�߫�]�.�v��z���@f�F�/���	�&������T�;�l�J2s�DlqeNk�C�q!#�0qD�e�T/8]2ꅘ�z!�\��ף6�o�LV�se�3f2�8"�����0��etSF&�Nc������D�ʿ4A�(�ki|����cˬ09d�a�gw���8��d%�5�XB�Si��@�|*;�#�<��?퍠]7�P���������<�lhdԺ���9��N�CU��V�L���CW�VWn-�Hӭ�ǉ��l�G巺x���\v��?������s&�����D��y�e8���]Y5��������.�vƠ�S��f��ϼe[5���o]&�^�"�����[��R/�쿶Z{>�S	�`�2�3\<��2���sD�-�GN��<��np���='�b� �|C�y�{�$�@h���0���^*r��O6G4���r�O q����ý�>�=�L\����=�8qT8��τ�����WX���g� ݏ=N\�%�3z�s܄i;��>�#���;�k�!/�w�}�A�3[�$������x虰�����������;�g>�0���;��3a:R6/��Ď�ߡGz�΋B��u�h�L\p�S�����BCτiD��-Tu���U���Tm��P��K��.~U�Zկڻ7���}ث�����PK   JrX �/��  �  /   images/25830125-c098-459c-a621-2bf82c8cd0ac.png�p��PNG

   IHDR   d      ٍ�h   	pHYs  70  70}�O3   tEXtSoftware www.inkscape.org��<  IDATx��X{lS��ݗ���8�Cp�&�������A4��Ү�¶�n+�j��6��P���J�K�
]K�Pي���At#��D�Bևh!�H���'1!/'v������|��kIu�5�D'��s��������[,Vt-	%� �｀�����T9��:�//������_R�@��~���U����4��0�1���2l���;ǎ������ t�`��^8%�F�Mi	,~A}F���-E���o�>����vy{����]S1���6(��|�D���w��X,H���c�9��<���E!����U�ա�u⨊V�ոf��D6!C�H���+�c��o [���Mζ�wn/�BOe��w@~�4��9������ymm-����!/�_�����:��e��jаS������R����O.crb�<�g	}�����\�����2	�QP,�e��˩	�U�}�#�^�ٔh����2o�iH`)�g��aHQ�+������������ٳff������g�M��瞻����BJ�tQƩwO��QyyK1���(�a	���B�`C����-�x������](}���G��!I���
E��]�+���.M0��E����
���AA�����@�x����Vp>���j�����pl(((�����(���V+JK�iM���Ca��p��<�Gn7ՒDSSS&Eɲ�P(�?vaY��r*+�UM��$D�!@@�^��hf���PL"��-/��2�W%�z�j
���l~.����\i+)#������Ԡ������t ''�����e�����	3s�� �H���dM�@� B�+�J��Ʌ�?�������(]^�ѱ0D�)R��t�_8 �l06F���U	D��*X�$ٚ����ϑ�
_dOّ��zW�Z�+--թPX�ژg�ԉ�D�l��LT�7��X��KJ�ĝ��+3�"V��,fc6 \����MΗΜ���$�i�AV�I�"�&��c����um��͵2X��ɤ����9H�	�����Do,K��� -����8=o/�f,E�8�t�
�Ud5d�������p���6�(ͅ�c�U�[x�� �ё�sС�� Ҁ\��),,$z�>��ظ���� �)��(N��3q�8�� ��vB�l���&h��x�?��y�0�O����A8�)�-j:C�(�C 2!�0������8�u����dQ�IC'?\��iHA��ʬ��ȫ��} �?��&cz�Ҽ��v�2�AGGǎ��J���<�H$ZW�X!)I�A�uH)3�l�t0���$����A�C,�sI.�r4��� {�%�^��@�\Y��ofZii���7:�Y�q�Kf������W&�+[���IC&�͈DɈs�H`glx~?��ټ�D]]�{�ȑ#o�i��׻6���x�����*޻�G�lR�x?�S��EW�>�#�2��6�>F���^���,V/��]�G9�fl�iSլ~:a;uF�Y�,\��6�ň�|�i!@�����S���7&�a]2<;��[D=�;�ʅ�n�L`E���{#8uɆ�?}c�~tvv��m��&��;w;���߾��B\iAHZ�N��[��E�L1����b>y��d�Ν�QL�c��sblRE4��X¼�*q���ŉ��c�[{3�;�<y�,�k֬1R�Kģ����=h�6C��/����eam?��c�w�MӥP0�������q|t�r8i��7�$��N�8af��%�⫇�m<���n�3;��^3�    IEND�B`�PK   }X�_B�   #  /   images/530fdb4e-21ab-4901-ad86-29119845d103.jpg�teT\��mC��Ҹ�Fmܽ�	4.	�N���.��K�7.��� !	$9����wǽ����ػ��Zs͹V�Q��H4 �  �v� ~� " �X��dd�$ddTT��44��T��44Ԕ�+5��������@M�"����+" @�$*)�/��/�����GDH"!��`bz������/������W��_�?��]�z �8�Q���N�$E�5 ��׈��[�?&6:�ޫC@Cb ��p01�����=)&9��%�����m����Whjz�4��wC�(XQ	ֈ�~�<s�^�Ǯlw���	�����ĺ�I�ޯ�q��@tL��H1��)X��S�0)m�B�E�XE�zQ[`��ƾ_� �,R )�`�g�j�%��;>�;ص�
0oSP�{�NV���S_�/�&�tCMk���UOj��P�!+4��z�_+��	��c����AӶڿhɃ:�+�o!x�Q!Ʊ�&�;�3U��͋$.��k�}������vl�~���·bl�� 50!0A}�觮t~J�#0%k��!�D*�P\pej)����3���FOuE�'�XԵ�T |����?9mP?~��׸3���tLƚ���ߟ�D8e�㴽/0VB�{���Rv���l���B�}�S��n��jyHdl�m� �����<j"�M���t�<v�u���R�*�bF�E3������H�t�0�CG� ���<L�yy�VV���ìXk��O�?�/��B��v�uW$�ɷ�|Bx/>�EůM��ڬߟ�<�+����Y�������u:��r?��e�"��d�o�B#�8@�i(�)�Z+�NDg���3KHg%�UKaK�$��x���R��VX�@��6���������P���R���]�����h�M�3;cch͗E_���.刦�L�������qڣ�@�m�[M�{.��h��֢OgB�g=��vB�K�A��6����J�����Q�q����r�l��QT흜klq��jsYf��ɩ�����F�OHa��¦Io�h��,���y6}h}�?b� ���D�[��W;5������i4=�)~S����;���(��ߣ��;����
��Q(���D0�)�"&}�w�2�Ϸ^��m�L�.�B"��'g���0�e�8�{�v�=N��lj����1r'ޭ7u�9_ЌQp�P���=�yҙ��S�x6\5�����)z}Hli������Ȫ�_�I�
�MR+���V�	K�+���
�)��a(�gr�9Ğ���F�D���� ��E�A����ߗ�X����pU�C�=K�U�R��&6@�Y����V�}��6%�_h�L����7������-`̌ �C<�5+�aO�^���,�L�����k ��by.�Qu�8g��:�8ি����:���=�gqp�����UQ�������7�?Qx�b=bSK��F$}��\��UV8����U�P"˼�a��]�:
�D�/5W�њ�ڷ�o唕�]z�^�]4��Y�n��d%�J����d��4�-~�r��,�E�"�8׏3=CQ��m���ߌ���6&1J6���@,�,��a���)	��P���� �����߲�����&��w��G��LW5aw-�@d�����U��"֚N��Ә�!(QU��̐| o����P{r��K-aܰ��)��c�U~��N���!��b}2�<T�,�ݩ���.ϐ!��ׂ�g/#�����TC��EȄ1h+S�X��WR���li�1��y(��x����j0���@D�j��&��\g�%�)��ڂ_a.�es\�y
�Y�C\����
��z�^Tȿ(�`A; N�e1x��Co�?��C ٷ�������#aD�E��3 WLxmF��s3c��ф_߼.S��5���@k�c���O�#s �0�m`��M��']fl�՚��<��{�{]�je|��iG�_�,������4OgN�۞�ڴpd�k�;�B���[v�� ��l%�汚����rvs֤����v�ǭQ@e�;��ǲ���,�oLThL��"��p��7�h�.ζj�3ZI��5�y�<��%?P8��R����$6Z�f�c��H"�̸U&tf�=��)Ƅj�R���F�-7�E��f�dй֕Q"2���9��G����i���CrG�R����=�����_�&��d'Z���
�$������c����*ݷ�U��c{�<"&S�Old�ր�^��-��^��G����TlEI��,#d��p�ǜ�]L�Kx����=Jй)!����|24��Y�t>։��?\h��~$�)��3��ϗU���nMS��bմr!�y5���1�!E$�@M�l�ǀ;q&�i��@q��>7���2$�`�qY�Pb��R�67���s8������i?�ѧ{����;���1Q,��Z8܎���[?1$� B0{.���yAw����%�t�3��J)��ګ��!BO�����%�o�c�R/��FG�Q��T�E�]<����WB���v�Q�2x�be��u�M�f{LK�h�-5j��[���p���0| ��9�D���OSy=�>{-�y�U}�N��&L9%�Jt�xX��|����6ۋ��)��D�"+G F���$�f�	!X�[�ᩭ9B5O5(脉X�m��`��jj^����Xt��ae�(4�̧��N�SH"Rj��G��l�"��pSŤ�����rc�H�,�	�rKǬ4�K�g��ڕ\�bui��k����aE���(�ƇJ:�ܮ��u��g�*g뚶��MeWU�&��+�b�\W�[��:@���w���%V�mM��L9�M"_F��M���
L(�>5N<iz�U�a-?\��X�����]6w��}��T�N.	1�ȣb�Y��D�(��N�+6J�	��Xz�,zb����t���ܮV/e�/�Di8�.��yw�p����<�z�h���3E����n�[Q[�����,͓_�M�+7�Ɔe���5m���vswъ�8��l�D����S��}�(�>7�V%8�͓�I�S�"$��GcV\�@Vi��U�{+�Y,:$\'���ɐR�dI�B���M�Md�΋�є1�,�<�5.��DU�~�_d ���R���H	����;��e�<�ˈ����t�k�jX�a�+�%�,Յ0�48��٬��{]��Tҳi������P������W�!Ji�az��G�q(L,li�5ދ�d��t���|m��q߽����)|(�P��|��^�$߻!G�z��y�d�ŻF�H�C��꤫*i��/g�9ڸ(Z'�c������C���km8&�!���$�Ѧ��֗)-wE�S��_ZQ�ɯ�M<k#�M�[�xv�$$-��s��j�>1U�p����)%����>�Wք ��ܵ�
���(��d�D�㒙��']��$,��:
���p9�L28���Ͼ�ys]�m^#Dx)����ʘ0�ܴ�qs��s�_|l
ۊ�������e�����Nmw������hJo�΅S'�����U�sHWJ eF�Z�i�iID����1./��Я��ysGC&���#�aq��w���E�j:��*����Z�^ ԙ�7R*���K�f��8 ͻh����^��0n�`��A��"�P�Ƌ	�m܈!��̮ZW���ζ0����m(&W��\���vC�1�.-��N�@�o]zg��J�+��_��VCv��yG![�z�Pچ�����*�z��p��YfM���
�d������|��唶�,/m�N�b��>+��q�%��T�BR�@u�N@N����'6<���N)�1�b���R��J$��_'Km��?i~�H��о�m�ʥ��,,0^P��I6*�1J���>���u����^P�t�ɟխ)����%(U3��]��63r�U��'*ah����^�f�1#��=xӤ�[?���4����b����y���E{T��0�K��I��6,(�#O����Nչ��t� {���疐��پ��`2�^1l+1Fe.�����n���Y�X��]x8/7�*"��_������b�A�O��֎���p�j)Né�ܶ�H� ����TM'��-]}���)�(wp�N,����@~$kg˔�����u0�櫊4�A�K~�T ��}K8"�,g�?����
�t�������2G�^*G��4�~u��w{-j����� R��c�!���70f%A'� Դ���ug(���3��ɲ\#��Ъ���:	۪,����ӥ+ͫ�b�%����wCs���O ~��6(V�[�ҴX�R�6��gR�d|���^ިGN=�e�E�5 Z�U�-��"��Ǩ��L)Fd95;��s<$?#-��g��G�������$���|�Q�wk�QU�"ba��1�b��0�>���&m|M17�{߯RX�><�M���&D�xn���5��I���w�=���T�'X���d�f�	f3�\8�����X�0'�;��8���zG/���X��"Y��~=[�5�1/O���N�\�9�? �l*��k�r��^�:�p" #H��^c�B'�9���}����"��ƭu�<r�]���=UH@�L`k��'�!YԬ�Vs	Ư 2w��W����/��D�S9��߭���^�C%�H�0�+�jy�
��rlП����.�[	0�(�"�y*j�ئԵ��i*���6�[<@+cr�+M����,H�"%��og��,\T��dB(��Xj ׉c"������n�#j71�]�����_ <�K���S�����o��\7��o.4���<��ҡ��^�D;c!�fb����4)4��� f�5�@��ɋ�D�M�h���NXQ�{��Gґh�k���V:�wSmY���r�g�	x|�`�� �6�y��u���@�ol=�į-�@�?�}�d�Ⱦ��౻#��,��˳��c�ʘ��q�-��?eI�sH���n ֠�� \����7��ɱ+��!Hh,ս�Js~�xHE�i��L|���KPQFҬ���۬�!����(k��&�V�g��g�~N̺�~�r�i�'�����Toy�g\LZ��*��"[�R�]�r9bIdZS���Zw+�b\�AK��ĸ����7�����I���-�28���A?�7�#�Zv���u�y����md�,GOԑ�.屏<ƽ}m��Jw;�
:De:YL���e��}�MX��j���k*
X�h�u�a #17���?�hm�%Xj4�����
y!���ͮ �LT�;B�!S�����C[�)rnO��	Vf#U*bM ����D��h^t�f�*��D�����)�	�C�Kf���p��s����M���.1n��J�#!͆~-����Ж���ic��%"w�,^�/pj�a^��n?{�j{�Y�_s���	B�Q��@F�@�s^����yb1U�B�=�HF�6��[�i�	Q5Q58���`���a�����&���i(�>;`3��Ht`C[���w�3���?��vT�lI�� k�b@�/�Ǎ[`o�x֢xj���Gh���{�咎{������)\B��҇��r�G��R�ˈ����n?�o���/3臖��]о���z\���A��t{y(��4;	hCP,ב�=l$���e�� ��I�t������b��B���R�b]49���Ѳ$�@6�f����}{Y�-;ӽ�=zg�r�wh���[(��u��H���le�	��yyU�uO#>��d���F>�Zҿ�:����V�_ t��/� �#��/d���|����� ؛"��wE�ߋ�9oƃOko=ߧ�.-�, ��7 ���τtxT
?9'���~ڒ���䏻���}�Ww���T�b�s�q��-j	��C��>�!��_��ys*t8�]^�_�O�\W*�i�ߍr@AC����W�깜��m��4w��벓!�8HuR'�������˼ĸ��F�����G��^G��AB��1�=�wh	��S�����r}]��(0��b��ԢeU����wLm.꿺q�/��[xJ5O�T��F۲���c6��Vt�6V���w���YlK,'�u�+���CU�p�h�-�������֌�z��Lt�d'������n�~����#�#ׄ��c���^�:7���|zմ1�$�՛%����0�t��d��<(5M5y�;rБ���yBl0�'Ie#��/�W�����{Џ���jD._x�~s�!O�6�*��h~6�p���_���:j�gl+���Tj�d��Z���KWv�u�;�~w�̌���(5�P�3���Dt�$/nZA>R���/;5��:���(5�w�����=p"�t�.�f�ol�⠜t�|u�f� �����L��Q�ql�g�2d.�P�j�~�uF-�\ov��S��J����̾Q��q�.m�FGg�E���Û�3�%o}���q/�������6(޼3��k{/���}M���y�p� !�}K�G�4�����%0�����}��i�?Ϻ��2
�h�gy�5"BYX"�ó(P�OG��嘽��&d%1��`�@�����U5#�e���@m�̽C���2bw3��/�d��q��J|��%�<�
�E��c�=1\֫����d:�l�_���ʰ�!Y��wzYS/��z��E�E$А,�KHg��d�����|��	�d&��c�,�Wc�R4{y�LFn/��Xk�4-y���ٶc��y.G��X���D~���HM���+>�O0�Z�Ҭ�(��Dx�_�p�?�����c��h���+��|���=U����{UI��
>��w*�w����攓�x8�ѽ��_) �˖�+�%��������]s\s�q��';�����Xؒ8��k�TqXTUj�qɔ�`�j�^ �7,z�������swu)��%�1�-�̀�V�N� YH9�B�oT+UK�V�V)���hhlG�/���AKq�-Ӛwۗ��+�����+(ރ+����b�P)��SE\���g�g-��x��?��ucZ5��]mOn��>�Q�{KA�:�|�ִE�\?}a55� ?�A���4(>	��D�Ƿ܌�x��${�,(}~���Gܻ��*����S�O�_*?�]|�i�cY4��=śSȂ� Y�ɖBj9��sC��`Q��@�� (,�/6l�]��� B��@�����J�����h@J�-.~��p�v�j���RxU;}:��=�3Q��dw�\����SXX��Ľ����B���R�`e�����ќ�(hsI�=���a�8.b�
�>*�u��~������4Zl��F6S�3(M����3��jϐY��)Z��eCE�Ow�ut8�~)�۱n��j��Q]$�BѦ����q��gȏ���
.;�;_[���T]�^��������i-�o�:-��H8FE��?�XX���.-	j������6�=�`���/����>��~�7��`���L8��ɕ�U�_"������5cTH�~�k�筂����}\$q1q$�Ix�<����
Iv�P���𯭸��:�->�����E0^��Lt�����V:��U�©|���PU����@0�yg�d�����tP�@��cOx�V�|}���$}�[��|���Q�,J^��N�(���!�����f�\v�%��C���ޓR�����drt0��@����7�����A�T�L�w:�BofO���}��g�)�]�	0gNF����	��yt�w4Nf?�Qm�F��/��aLf��|��y\�C�]`��᳎Ԉ��.�j��{l�����}��6�*�O!���kw���Ge�[�/�����|��S�-�w�6�?�?��w���@C�85�u�����F��L�N�^`Z���`�w��2Ǐ�l����-�	V�6��A1٦���o	_�F���Q�ˊ���O�v��6x���р*Y�*��Gi��'knYv\x���Q̸ƫͯ,�Q:����[�o�n�г!;+5�syK��@���w�idd��n���b$��³|���d��g�t����(�t��2C�=X K'�Vċ1�[�"V'D�.oQ������B/}�����5"�,����uN������5�������Lm�ẘx�Nd���I\[��(�L.I����s�*�"ЋXI�"b�"b���\���6�`�Urhs֤��wA�:��v��U<B\!(wzU�� �� �m���*��{�x���n��;�]�����2�MKF���� PK   }Xv��^}%  �)  /   images/b7b52948-3c4e-4eaa-8c83-bc90923fe796.jpg�zTSݶ��(��J���TQP��JQ��
J�.HED��"�A�� - *�K轅�CH��_��;��OF�H��{�9��{��FB&OG5U5T** ��� 2
x	03b<�����x����Q.����GϜ<u���9A����_V�"|QV������,T��M�+Z�5�un�T�:D��t����'/��>s����M �!�ا�:P�QѰQ�[�2)�~]��5-=�.�Q�������������ė��e�;vV\����C�s.�Q���K?s������5�����S�\�/
	_������v㦊�������{�F�&�V��X��ڹ=s�x����2�U��7��1�q�	��2��g�����TV^QYU]S����֎������?084<2:=3;7��������������P4T\������������*��?��ҝ�?�������9��C��Q�������x���t�����͟�~)��	
��R���?��G��4T��ѰP`����{0�D2���m@�7���]u��`̭�B�(>A��� �[Vz�i8W�=�Tt���L�1�mN=�jHC���!��[�p�F��/��Tه�U�X%�1��a܇�>����p�C��+�>_��j<�=��^�����&2 �����Xj��A�
�3f��d5
yb�zK����I
��hܱ� 5?U��ϳ�u��w��% &nоQ`�����D��J�4g^?խ�krɽ�H����]�暃Zo)��9C��vtZi������`��0fc�ь��u9㗵l ���7�����s����գ͕�+^�1,�[��b �o4@�,�`E�a!��uʝ���kL�.E�?D\��J�2�VK[���'���]z�����BF���	�c2���oA<Ѯ�z��uImJ���i/��Ѽo��!I��y��a��Zl�Ъ�ᐖ��uZ��|���a4v�f�ߪm�W�#����+k��D�O�g0T�0�@�I�g\}CȜ�Ͱ�
� ��������X�4Nf�7��R�M�hcOKK�OH�zQ������v�[���b��U3�p�#�y���E.�\����^w����]mBˈFCr�������`n�i�R"�feWa��
L�Y��/#��Ծ��S�0-�75�~j�=�nq
J��(/����@4��k�x ��ǘE!�����}��B�3o*Ǽ��'�S,sj����\lB���_Q>��9棗o>|�h�u҅u�����[����,J�,f_(*Pss���~�������Y�Ӟ�|
_$�hY�Z�l1�Q6X:��dc���(��&^�o|��;iM��*�if� ���f�p�f/ڶ�A̖�C��)��t��n@:��t@�4���q)�H��7ɿV�Dͺ�E:�J���ɀ���������Bl0Y��x���M `�T#MJ��`���]�8
�[)�e���M~�v�����X��~U>T�O��j��o�n�&�!B��(�1g#!x�A��VA�������&��J�rq���-꒾�z��TG�;^)3�_[�����( m�"ٽ|ܺ���#��R�~K�R_��(�e,�8�Q+^Q�Q����`����3s�M��,9R�u���^M��E���*��u<`���������o����m�mj�b-��+*=��� �뾆��<�<{�@��G���[�aal����W�-���-���!����^2Ь>�C������ d��a�q����	�`�o4d�\�٨yr��A���*5��3P��h'�@	�C2pٌ��,�)Ƴy�>B����Ӂ+Pu=U�[U=��4��٣�����:,�8$Fa�hC6���TϜ��Y�Ao_4x�''�._����zTA��)��\�Geo�ܱêcgo���FR�ʔ����x�Xb��ΐ.ݿ�'�+gl���$8�cU�lOd�Й���s9��Z������E}�c��tF�7O�������x]���H$O?(M��Or'>����LCH�"9A_<4Dѕ�w�.���ߝ�:0� �fp�3e�)�Sم���ߌH7�X��w�~-��Kg�V��p���̬9�y���cI���>V���~�=U�슪2�>i��*���"��Ǜ�W鍢VV�4�-^�нi����2��Hg�����"l��;��*���w���ۺ7*٣�5�;�>��J��xN�<���:��s8�1dзΩ��0�mK�	�t�x�e��jŏ��4���%�Ĵ3�CK� yJF���:bv�W��z���U���T��O�ww�U�e+�}i����
/�\v��4G����F!@���M	�C{�N	��X˺�1�q(�p��{(�lRr�Z�L�-��UҎ�v�J�[8c*�˖L:��Z�p��j��Ju�[F�\[� V�w<��LL�,��Qa�M�Pak�6��)�ʼ�8��қ�oYjz����9{�^'}��s6���\ץ����j�Y9Y��U=�og?�N�rt7TO-~P���K�A�}�����u�m���$t��+$�BS�]�)�b�A�U"n����R.)���D����N�j(^aa�+k�J����'���ߦ�2~M@����@������{�͌E�'���#�"���Y����NH�r�.��,��������*���7sN�ŕ��QߗI��ѯv�����d�	�Rf�,d�<�p�KąR�S�֏i�4��h�U��h?��R��x-�8*t����s��,U�/�n���l�x[{�\��oyfȀ��u�Է��ru��䘸������d_��z���j���G_(���v��Q�l쮠�x���G�N�{�1�Y��Ƌ%���k_�Z�����T/�\��Y�[�ِ�r1.�5���0�;�6����v��QӷR���;��Sl�C��K�_#��"�?����}u��;�2�q�1��yw#K2�N!q,{�]�TY��|�pC9�`�S��C�쮋���>�w�.��<V'j��pVI��]��X{Htil�;�3pY�����VW�CV VS9�L7��h�ʕ�Zr��a��K��@~W>��R(����;��y*��/�ѐ<HT8t� ���ge��|{�^6+���1�"�ђ���w #_�� ;e��2��恦� �=��+>��I%�͌�_�|�����ؿ�z�m� �c�:�
�����24�N�X�$���h�}�ݲh��>;-�M2�ū��3/@�9��`���Ն׿��`��ꙿ!����d aM���8��iW�!��جO�
�K��J�=]�4^C�
���b�0�_����L
v���m���Y�z#�Y��9f��e0A);�۰&C��(v�pme/b���ٲC��n��ն��]n-�C�O�����_��E8�D]�d7y��6'~�Ee&����~gqB��F����`�dc��,q���G�,C@������z�ڧ�d�o�_��<��l�;䴾g�F�FE�Uu��Ă�a#g���^Y=���5܈y�;��:�w�������g�Y�,��z�ڙ/��W��Z}���t���&*'�#��V��|��(��r�� �	
�e�� ip�¶��od��6S��˘5Х�Մ�5sD��@UNbxv[^��~Z�_Z��ٜ��'�c�Z��<�I��Űh�����E|'��ݷx<$��!q�	9�S$tb�W'0�����>+GH��'ӹ����tUO_O )O��C�nG2|9&0��A�~��.]:�}���{�Wa����������/,n�W�����
ߺ�gE_��B*�H0����P�6[���{��n���uQ�*��
k{�hZ�Qh5���'�J y�!�v��f�J��8���b��"�l���"h�f�AW�b\�
��md��)�s����:�<� Ch��֐�U��$�!�者y�͸G�)֥g�z�J�L�:�j�&�lyLP�zq���ca�~�%�W�Fm���1�~��9S%g���V�q��F����c��^��X���T&e�ڑ��՞t���_s�o�-��I�u��"���ضy3��GZ�k��H�+9�wl3S���?j\�v��T^���@ً(��d�*ݍ�M�{��9c��^w6?.>��,�x��g&���$Q�9d�c�o�Þ��gɼ:�;j~s��#��r�2�h��ngF ���G �X:V���c$����֜Pw��k�b�\�jjX�r��S�[+��o�M �se�رk�4�����ڈ�2`G�z�e��
9W3���}���x;��#�pYe����3F@p�H;ج5Ս�JE̷�E��w���gB���T���t��𡏖��a�����t�)jo\���5̕�'::n�,�Xt3��9�k�������c9i�Ë%2�eJ̦?�����N^��|���>�TX`?�� 9��t�.4�����m��o������&�׈������"��V���xǹׯ��\�N)@�Z��!�C�3�%!]�h�,ݯ[���mO9X>�ř��Юm�n	���8�;��+��!B^�*�sF�)���>%zyM��c���2�_�G���na9P`U�y�j��������)�J����@y��y�}��Ɖ���g���Ow~	���G\�;u�'�+ӟ�8#y�V0�:��5;�y [#�+/�-�JhW$Ĥ���Q2E{8����Z�4a;���J�o�z�W���I�ևc[m&����G.W1��,��a�8C��k=��bR�.�)�p�Jw�$q.�o1a�nY��L\�#��-Bw���������v�`���սϝq{�s�,�mj�ɘ��QI�V�ԍ����]ν�xtƷ�����5���/D�k$�27f���*�X���o:+;ɶ8�𸠍$�.%Y%���[O��F^T^�dd��WW1,*
G��-y=���â@��ϩ^�%�tri{̌0�N�)�Sf�����Z�7�f�n.3�����WZ�^1��{OA�åo���To�U�~'�m�:2�D���!Sr>㪏k���
i�i�n8��=xf�dQu
3�^�1lbdF���߳G(Ι}ğU='��I��ftuf�q~v�AoF��<6�<R��>�:WpF��Q�����$nr��b�U�ח˴i
J�b��وY	�+��W¿\�9�2|PcjS)��}�i+��_�E���E��N����y�>Ժ��1�%v=&7x��vs�g��.�E���-H�n��8D���804z`����#���D.���D����F��j+�kX��[�x۽�
�\wD�Xƞ����g<1�ׂ&9����U�ow�>]u��r}��[KL�Z{ݳ��J��Yj�w
���e&��9^�%�ը���W�A�|�J] 4D##3E��Y�ğG6`�}v�ee���I��}�ߵ�rU!��@/��Jh�A��KT^}����VdgZ���b5M�BX��R�`�d��R����u�nr��
�i!
v���4�#�݄��L�V��,D&�^;�D��MU���t�K��ƹy��4 %�d���DS:s&�;�F:�z��{��N8���tS�^/{\�B�|�)�$���{�����|Z�Po]�҆���J������_¿DĭDN�X,mjO��N�5�D:u���>N�Lք��Bl�N�9d9�4V���)��g9�F��e�W�p����tx%$���7�h|�Dx�|�~]|1�n}ԍ6��ׯOT[P��Iy0L���F/wۻߟ�7�ҥ7t� ��Vd���:�䣉J����?�U���թP���O�]��k�m� �ޮ
�
+��(�V���s�S���[��X��K�t�ۉ6Bc��j���A!��Ƕ���V+к���Y�΄�ƲNʮ�����m`���{O�ȸ"KQ�����ǉj�$��z���HĘ5qE�\�؛�8���y���۽�z�ȓ�4�{{߬<��*���_�{%�3'UΓ&�!�4�	�R����c-א�PL����m%J�_���~yKm$b4��;z��1��U�;��[K�#'����y���~�A;����	�hA�0�kD���O�'�Q���P[u�;+9/���u�w[�M����?���>�(�����z��:8H������N�e4'���� �َ����}�-��`�,���X��V�L�hA�l�צj4Ϩ�d�iH̏��s� $Hw�>�f��L����+�����D:�:S�&�����.4
��.��糥$h���g�6s�4���T�������e�C����at�4b�Vq<��(����ͻ�:�z�}�<V��N�6����\?��똎:���pOsg�ʖ�,��Y&	� ���Pc5և�J�Id6H�GA"Ӂ ����9�P��~���K`p"	���y�@��Z�2.@R� w��DZC����3,n��&20S�}}�ަi�(?���]Q�W���@Hj����@s� �8�E�w"����j�	#��2�փ���Ϛ� �m3�;^��k�����:�K	GRc���H��Z����l�ǈ,
��M�]2&����2��)X��pAT��仆����g>�qAe8�����M��W`��@�پi����[�1?��x@�M�[��(NgG�&�5h��%�M�?���8O�3�I�iV��n4�|z.Re^Dl�Y}κ�ծ�wr~��������y|	n����<l����ԙ��LMf�a���jՔ=�WT�K�e�I\b�`���1W��0���}���žv�������7�fO;%	I
q�RݑϞc�1�EV�N\3uL��t~��iNl�V���K%�`
�5�غq]�b\ 1C���4CsB�������� T��.=��R��hV��}���X������c;�U�W����[�,��J�ݪD���uh��/~�ʡR�ml�zKZl�z�*�ۺ7���}v�"'����ٗ��N�+��|�hT�l��Lw6��SB��}�e��D�!yK�����{&����_���:I����8l�,�bl8�g���qfxy��W��� ~\�ޗ_�tL-6'�*Mi�Έ��Pfd �=;�')�,X���N����4.»� ���Ǘ5�n��H�ǆ"���n��qS1'�f����U��T󂋴��r��RZN+J1?������l�;0-�|S���t��ݬ����+q�_�$�狜���c��U��%�p�%f�#f>c�����-`��2��{P�37�h�ؽc��ر�
yX{a����	���d2p�l�8�M��?�g�OLt-��]�v`NM���X�uW0��5;	�d�.ɽtZ[�����{�ﰰ�NE\��3�ڒ�Z�&n�����\_�j�To�:8cF�-�2�x%��bf�Ϙ���tv2���{R��"Nn��mE�4:���~ك��on
�J�O��>TBf�$B��|"���;E�a�n.|��(��-z��Z��Q���v�p����7_�R3�2���E,f?�|HInpO�ڰtq�a�+c6O�6yQ�"�mJ�6��uqؐ-v�W}$�iB0d����*���nY-�b���Ff�I��1�s��Aؖ���μ�`��� %�q��?�������'��O�d��#9|�	Z�E��v�����E�9��_H��؋ ����B���$eچ��,R����ɟ�?l���W�A�.ʰJR�~�ǐ����N�	�s?�p�֢4E�ߩc�K�Wy��m�y8գ��������N�-\Hę���
��I�'7JTS�'��9���{�����b��<�>9�P�f�_�$n��|U����P2P��AR��U�wSd����	��z}�l��R4)h8�$\��t���.]�:S��-W�uz[#�Ψ~�y��<;���^빌<h�����$:�c�8����I�nQ�4�^��t�V��1��[A�7����A�Vz�}5�0W���=��,G9���-}}������020?D�#�@(Ͳ� >�D���~����?d�zC�!P��O|
��&=��`�ؽj�C:;D��%����+�n<A����Y7|��C�V�\y���5��m[��K�����t�gk�gk��M�tE��0c������N�3��癱y��6����5�Hm���G1��bjT�r'g,7߈4�9���M2�,zKw���j0��?���.���.�^�hù3���:QIӈ�)�
+��E��1�*��1M�h���)2�[���iqE��OЮ~e��X�"�6%1˓;��}2�:�2��\F���Ug!'���Ta����R=^��K�T�!?���"d�s�7\�����ek藭�?�)��m#5@J���_�\������i�w��
ptc1���lx�O;Gص��:���Ҽ�
^S��s�$h��ͺ9`�~��"�P
 >ѵ��]xދ�BĿ+0$�a/�W��L�-�N�!�K��b3�E:�+GJ������/7���]����x�j��k�؂ք��پM�?z�O���?F�/AЋ�7����.�^1����x���b�<�x�i��VU�R�r9W ���[ǔeM ��������*��,jm���Rv���V��ϵh�����z�>{��s�����[E��
:c�Bn�7v$�;P�8o���
u(v��%��֔��Wt5�*��;2�Y��I�;�s��63�U��Z�&v�mL�递�|)k� ��ԋXz`A��!�~�1y������D��o�R�l@�gw��Š ����#�@�T�{rI�S~���t�O(�!m�� &o���>CI�j	�Dq��(����g���|������!���N\�+�D9�O�D;��2��%����"}�Y-+r�+�p��������1{n���P�8�����o$?�V����t���J�{���H�uq�>x`k�s�	�$]�͎e��$�⿃����o\_d�ܝ*����м���i-�������*tz拠�_�9#�/3�_%�7�5�g���_��eɔ:Oq.k���/��{��fCįA��׭���m�������~���1���z���Cl�|g�#�}��_���ڞ�_]�2�eH<�L�%�p��އ�f��I;��
u{������{��MIy#���g|���,��g�%`���O�w�<�,�-$t����Qn�:<�3SE�)�>IY�����Tw﫽9/Xg����B�Ǫ��"���%MLZÁ��Y�2��N��KUMN�w���K���s���.��B�r1i�x���]J}��.�QW��M5	�Q��ӼR��"싐`��f���;z׃3�C!�t��3C���T��챷�ڼ��?����4��T؁����23�!R	����Ut�������x鄎�-jl֙��}�0��|v���Y�cI�7V[Ur_=?�Y��!��q&���e�"kP��A�乏��!�_���ީ������G�PK   �}X$7h�!  �!  /   images/c6364832-c854-438f-b38b-75bf2a0cd33f.png�!މPNG

   IHDR   d   G   ����   	pHYs  �  ��+  !�IDATx��}	�g��UYwuuU�Q}��P��ò�[�c3> ��L�L0��%v �`� &�{�e�X�;,`X0�c{| �u_�:�Շ�w�}WV����է���f��������������T,��~*,���t�4]М�k}��%��n �-ȡ(�a 5n;*�t����I��p۬�4(�-\mPh �����	+�~'�oQPNľ�i�xcx���Ώo�ƽ]�hvP�i �BQ�vBI�M�O�os[��ǣG��Z��):���H�Wj1
�&�&y�G�P����
l�]�!��kjW�v�!⒥vVjg�/9j�c.;�S��8����������Z�!��Z�r�Cn���]�(�v)��dE�c$ wQ�e]C��p:�X&��ܟb���g�ѳg���ƪ=7�vp�"Yj�͛���4��2�ES��t���#�bzj�u�PU��F�q9�ZU�h8�d*���F
����6X�ǋɉq4��L&O��pX�V������ ��)d2��7 ��c��U���r	>&@e�譼�l��Oc��;����u���F���N��?3����&\nL��C�����!��#	����MG�[�J �ӓ�SZۺpr��H�?E]��e1�Jz��4�,X����n��>�~:��~�K�"���~�z��g�P��Fs��� �ɑ����,l���CMu���MN!�&�"��bdl���̂������ëZ1�A�u445#G�G�g(�NL"TgEU��D*���I�Q���(*�T���pvzfi:�]K�P�6��F��'\��kUĉ�����������D�����4�����>�������sb�b���ghc�&�2�[��_�gn_U�	�-����/�J`�e!s5�w/��6�MiW��������9��V�}E(Ni[o5�vˎ�R$���������Ϧˊ]{��,�S���'X�@M-��ד頾��m;wR3����]]�kE8HJw�|Xu��6L�2�����9��2.zf����ց���Ј&��I W^ú���zNim��Qơ��7�$��Q�Vw��K�x�+aH�/��D�ӊF�!��׃�-f�^�����6�0�
�Ȟ�T�i��b�#��]{����ؠ>�^ ��yltR:���������TN��Ͱ�%V�l������D}b�^ ��P�!E�?I��٭"<S9�G��4��Ժ�ই��E���*8cYN:_A�K8S���������	�T�@8����Z�FLq���fY������̣�e�,�8�����+e𙭝0�a�� Ǿ���*Ih��!b���΋VX�T-���܁�;3q�ܕȸ|�OC'�W�"@��\�7����8hGM����?u��c�L���at��X�ž�!��u蟎b8G[�_��|4��σ�j�ʹ�r׭n� ��DWc�^������Xa���&���i��n�h&b��������p��)2Y��n���(��0ZCU������R�St~(G�cS|t6V#20
�|-ɲ�&��޷wv��K'�\��-���/"569/Wu��yr��ܻ6`Cc-~�IK�tQ����a�������Q�`��8�?۹��n��p��ÉuV�omD�ߋ�Q���y1��� ��"i�A~�D��"���z�H��Ɉ氆��۸�p8���ؗ��@i!JRʖ A~������훘�1��EX&#H�r��
��9'�#�]K�3u��dV��M�B�U�d�tznT�gת:��;���_CX�;~����UȒ�fHz�^?Ԯ �������&���!	{�yZL��Ldɜ�p) K���5֒��[%3�����;G>�FDIҀM�SD��``��찘���!����vS������/s�� p�:Gj�'P�/�&�M��i7�nchb�f�@)G�Dc�Z$�ŋg����I�Tx�:X��3G��O���
4��&ȖO�T�J�w�ā�29�R�f!O���T��pD�3���H
llO��g���J����A�|��Y,��q�LG�$5AB½k	���e�>6!�E�p�(����Dd38�~�)������89|E>�%!a3�-1�+K2䏫S8�y`3����h0i�
=��*ND�񲽎.Ē%FL%��$�f0��y=�U:pa<%���'F��T����Q"3�0d`�/Αy1JQй���Re�G3��q��_��x#fHһPi��3׍��Hr/E��v��}�E�H_�}g�_��H4�
�7���^��&�7�/|�3�r:�����Q�mU�R���J7�F5|;��hO�8'.R�މ�t�U��6���cf�.�Fj=�'��
}�"CIg<���k��i��XZ8M��7�	|90_{�Y&�R��kT��X���cqS�8�`Ma���f��%F�)
�@b��͎��o&~���^��b}R)�~�����i3��[Ŗe�d�6{��2wŹ:?̜6aP�HD����Z����8�:�*�Đ� MQV�� =݃H�zd�������)�T��i���
���0m�n�m�ߪ�yE��ܰ��R��H����,6Al"��EÊ��!��33x���}g�Ŧ�}�!>����^��߿��`������f�q��9��@w���lz7]#g5s�����M&*�)�e13H*�>BG���)��ό\Y����m铲�L�M|�Z67L���c�3��i3���%0[��^[W����3����;���T����.m،qnB�1J݂����&Sf���.�A�b��� �HI��?,�q<�f�M��#�j���6F��$�	_�4�N���_&ЅXɳ%�d�&����KOh6�ia�3OJ>�$if|G<�t�%y�|�d��2��Y%fVy\r�	X�r�(0�����'�e�)K�+��Vg1��o��;RrZW��2ODy�3�¸!��
��Y��̌:��a
(�9�ϻף"�	��_<�,�;O�.�:,�;���={$�LPd��g��[��_O���ޛqφ�T����'��S�"���6Y�_�f�:��x�#V���9��
�6��O��i�_�TpqYy�J��gfwi)ib�T�n7��8�**)y�![�#����(��9�է��k����������ַ�k��6������|O~�����>�<N�Na1��o�h����I�vܷ�/�_ ).P�8�5uAѲ�(9�g�͉a���7v� �Ç����s��5A�����z{°��
�;N�G�+n��+2�W�,�y[�����6&��{_L�*k��g�p����?�߱A�;���Dߵ�_y�5��F�v9(b�r����V�{w�7�w<�OߺYL3�����%ʸ�.'��Ղ��g��˓��f(�v�QM�S�mg�r�;�S✍33Ù��y�1�Ḛ��������a>��w��|��Ib���~���q�??&����;�Dy�NSҹ}U�� 9?!�R����&�Vv�ϝ�~����!��5�)'%��p�n1W�f9�˄t���;���g��`&��.:XӾ�g�,��O`)e��&��9$-w�5b߹Q|���bj�8އJr�~:"�񼝋r	6�����lN��a|����>1�E�*���}��"�eq+O�q��eO�����T�t��4���@�L&�a''j��LL�w_;���s�H�ӽ�"�~/~��$0����>x�����ɡ�����o���i
8*ȇ���,��5�w��sz<�f�O�~6i��L~���)�oG�bKkz��1�|�Qr��n��l
�N;O_5��={:����	3"Q�kM67Ւs�P���ϒ�'v���i�E������I]f[9�������XC��~�%{��Ħ���������\�W�>�g��)\Of��������L���������DX�88`����Z��x��1ay"��hR��I��>�έ���-��()��ǑD@�ߤ)bc�V0�8�i:6ӱ���WOCs:��o��M�����H�9�KĲ���K�$>zC'�m�R�x� ��et�cPR�D؟���Na+K��<�~r��0�CZ��_�S=��]2M��C�(2�EI�����'�%�[]���5V��7J�������sp��Ϯ��m��ZC���FN�tƇ��G�Ã��g���׷��J������ꁫj����aUE[f�(7����Ȕ��(U��}�~�L�a���������x����)�1~��*]v�b6L�C��?8.����&�;ֵ���\6��'��j�y��(�0�Q���B�"_��,}���1�e��O�|����{���� �0-d�9�� �:�Y���DZ�ſ�;�H�\�����0�P���3�s��}�u;�r�whxS�Y�3s֞����	?�
�g1����3�f�,�2b3��9;�����\�(���KG9�\�)/�R�"�&���v�!��N&kϝ<�#S� x�-�cUx��,����|t��qe$͉K&
;y�����7��P�1TY����_��?�c'��O�V�U-�G�lUf�후1f��7�/;DժcY``���RT	c=�kJ77����?8���LV�M�Uʢ9lu�VL��U��*��('v���+��1c���1<�8@��a��t��m�5E��*j�+K3Ư/�����W�%��"�q��hּ^
{�뛜i_{��sU�R�S�g����ǥ�i�J(����� �,/e��V�S�����!�ݨ�o�
��Sc���4��{&�%�%�뫊�j�Y_�7`��0���~�"�.6X`
f�,�]�av���	��<��N�a)de��%�	]
l�U�N�4-U6Y�W�MNY(a{z�a4��OMƳM�e��_z@es��@!��@&P�8C���IWxkjq����_B�߉���D�u�^$�9�ۄp�*���s�h���ܗ�?0rA����ZWZ�H�"��3SQس)xm�+01�&�VDc�#�t��W)KGY�?Ȝ� ����(��0���ݕ�ȫ�u�|�~�"r��j6`K3Ģ(ט�� I�j�n����d��J>�`��n �B�������A��	ԫY���	/�>�E��7�`x`��Q�<U��VC��g��C�Hd4:~�\�Gjs�g^M�� ��5�����"'�[�y+G+�/P��J�!�xE�q�D���6 3%O�F�3�XW��32;���Sqb�&�W_c��<�hXuEJY,<����y�r�!o5pt��44��x�@�����]A���q�D<x�d�-`���ባg�/R�ѵʂ�>���C�ష��`������5��Mp�s�o�!�L'���(-��5X�)���~����S��*��?g��BqW �鋬����+b�;�w
�fL��czP��a�e(�p�4����h/Nf���K޲�w0���^��p��&��(��U�A�r�HF���D�S��	�v�9s��J3��wbP���cE�y�v��>�f��%*�	��"2bN��L�����hЋyٵ�!&8�S�nyg�$l�y�X�2s��_��*�*Ic�;��O5;PW�ď�
x9\���+�_^�E�3�ك�D߯|DKn��etD�:��j��~��3d�eAe���ɂT��J
�5�,��f�t^�7�sd9�ȥy���J٨��&;Bd�/`_�L�5�\6,�!���"��)��y�3)r\�A	(��ȼe9Hi���Ey�-�>D_��Wd�d�P�@�e╡�RIC��{.e�M֬�l�nW޲n�ˇ�����H(9����iooG?�<�_�#�5+%0ʢ�H��:��t�>��I(���//�'"&��TS����������*?.'�V-Hk���x}'5���y�T/k.]����֟;�h�.?R���^�9ӊ��ͱ�#��=pU+nڸN
�x���8���K���P)����E[[vw�¾�!�9݇�@��a�;�)���f�[,ڮw�z��
`U�Q��-�y��RE���̓�u����&pv?~����GQ][+�b��Ə~�#|㕽��l�06��g>�lٶ�͎O��G��K�����68�,���,ʐ�7"�H�)�סZ'��Hj^ۥ���V͙wfu��ަ
����B�q �PY]�O�٧����'�R��/��ؼ}�T��
1eˮ�x��
���p*PK���wf�)â9r�:::f�s8�L��D�Uu.*�#.2)���ҥ:�������e[��~���}����m؄M7�(eYg�#�͠���ݲ'��&C}���[,�� ��t%�K��`)��w�L;lW&_&��/$/�yn����aF3f3���5d��;;.Q+DGWW��=s��L+��1d����rŋ[0�0�b_	��)
-�z�p��5���bb��9߹�z���D
(3,�~������|��\�@�bL����R�*�%�xAx�	��}���r�̮�S���^8;,E�̂2����|ny�|(��]��(�Y�
����}��$:M������*:�8ݾ�-���a���Lb�G�Q9|���=s(���NI���G҈ݶ�c!Q3�4^�u./){x[3�Ul������q���9���2Q���Uu�g�9��p�����0���C��Ɍ�]���0Sjp,���r�j��H�pr�gNJ����]�]�MF�ۿ��fHYfCAY�u쟿�u|�k_C$���0JUB!��@���Y<���bt|�d��֥��v���B��ٚƛ;�LDG1���$t�E�/�]-XᔭmRN6�Ɛ�ʮ,���-.Zz�պx�i�D�P8.�)�����'�A��q�cޟ/����l���cH�"�C�_�iQ\s�vD�)�ȡONO#�����p��Ĥ�v5����O"�JK�v��6��Dcc#��uT�r~&6�&<K'K��|�Օr���XJɤ`��2�At���|�R�ᩞ��E X�yK�l�[��ZޟX,�JD.N0U� g�Lv򲉒efŽ��Ic����N��鸑��\1���7�����d\��l�_Y�x۶�KE�\Wᒍ@}���p���ۏ��fX[6H�SA���և�SIL��M� �]qU:~v�t+K��$Ō�ON�Z����i:j��睷�q;� :#'Vs��c�Ke���#�d.��ppi?.��1���
`�|L�4��?0S��vz�v�7�R���.r����?C3��&�sr�!��^u�L?.E�C���y"�b1OYj� M�ʾev$�5�%?1��q8���&�����3s��'F�?Ra��:�/�I5_)��G䊆<�,ȩ�OFxH�:k���YE�a$T�X��&d+?�`�Of1_�a���ʏW�$�� |\7���|H������h
Vs�o��B� ���H�^�ұ����z̳�2���j�*�l��A��O��X\�X��YԸR#�Ҙ���S)�x(fy�ym8
)8su���I��Ǣ\N#�b�p�5�>r~H�tr(��8~�"�t�s���#�%A�0�	25�|��'Ϝ�����Y�d�5$���z���35��p�!6̈́#L��S�BOdq�d�
u���ӲAǫ���IL�I}����ǩ˿�t!�T��l*�*��v؛:68[��31���	?A�}�D��s�B��B�{�i�m'�������B:����)\�!�N���#)U��G�@s}O��|.�Օ~1s�x�n��Nj���e�,2��}>��}7R��<�f�U�^����H}I%��x�bw ��I?��*%$ϤS訬㯠h����J&Q$f��6��u���?#�|��[�!�<dl}/�w���b!�a���zq���dR�kJYp���YImy(g!�ǎ�su%�NP8/���-[��_�9��[���If��`�#���Ν;)�Ȣ�p\w�u� SvapP"�M�6!FAƉǱm��9&�5}z|#��c���8z�� �i��_L$O;MG#��b玝b�O�<���fT�z00:�����m�d-_":ݯ�uw�!�������t��:� Y���w/�4����]	"�ljS�}�fю"����mb�y������ۥ�-�=ߴa���		�Ch�J��;�m�v����5�;I�,bf�>�ھMp�RKc��ċ�I�wn�j��֮�܅���ڶM�E��o�qԞ�����͍(^���23$)�?h~X�s�bb�?����#F�,��_.�ʸ��P�V�-E��U�|����/N��Q�C\�����W��)yk�����[�߽�9��h�@4����fJE��YDp�g�]��Sw���n�m�F����a��7!�3d�_揂q���޸~���M�I��)�G�2�_n���"S����,1��d%�³�����1� S���    IEND�B`�PK   JrXPD> �  ��  /   images/ee20a1cf-a7e8-45b4-af39-6cac45e8073d.pngl�TT_�>Jw)
JK# �%!0� �� !݃����"�C
H7H�t��0��u������`���}����>���L���11@YA���u�EF<�������_��M�����<u\m=},�m�|||^8�8yXY�ټpu�˄JR��1�d��f�����f#a��;~ʅ�=X��ß�3�|���	�ɭ�S@[բYq�%̩j���n ����9JO��ك�ek�Rf�q��;x�\�s/Ǒ�,����^1��y�*S���q�*�pˏ� �������[n]��Y��:p���׭uMA+�$f���'����������7�"k�e
��t�d3���X/��[� O5l:�{4�3��Ը+�f��^1��/T{ݴ7d8��Nuh Z������K{�����L��� J|�uB��ӻ��p��4�%�)�*J��,��6�<*���(<�η��[XX���.��i�D:�2@���A-P��^3�a���x��z �$�Ha"Lj�,|��#���纣���� b}?b���h�\C��ʿc1�2���6KO��S����R��r���c`����	m���f���i���ézL�_^��"e�@��qjel@�A��VT˷���'�\�|��g>�~j���d0sI{��ix�_���@�Z殝?�������y�n��G�L��RZ�䋰����|yz�x<���q(�4ȹ��.�<B���#Kf�� +�y��r��8i��tϱ9~JPȺ3c;
�\*�A��&�m��(��~x���لfN�P����d
!<��ֿw�U@D��!���/$X�GmM_n�ſ$S�{�p�J�g*�M5�\���s]��.i��/��k��_�&=�%�B������F�D��wt���yY}V����J����Bo��$q�v�9+�
c(ɘh����FRY�Gh�X��`����{ȚA�/_ 
�ϔ�yщ����:�f���s��'n�9����N���yڿ�ھ�wv ;��Ӿ}c|�v������T�u�$�-nr�r����<���!�4�Ď�O
��_J��](�2��]��Y��7��6��=nm̅�ƫg)\�=�~�@G'��������V������c���������Xh�zo��
Gre:;�[<[�Y:� ��좎�B��W_�]��]pP�����ln<~t�;��Ā������43�}�bPڢ�Г���|�����G��Y���/"o���fm���Ph���y� n���̛��NɧM_7�־�G!i>����6�2rK�0|O�6X�RFq�B-��h8�,��
,Y4��W����j|�O���:=u,�yC�v8_��*Ck��G!�c=��8 ��6�$������$zC챠�$����h0,Y-є�o��ʧ+��s�H�j8��\��3��_㱫Ax�}�K-rF����_������K$�>��
��o�l�T���a35�����ʷ���Xj���D�͉�F���%���vZǝ���c��l\��ݿ���/T�k�ΝTWWW�s$C(&�Ŗt���)�������
	MNO��������4������zz{�23U���!�ҡ7��*�����F��q��r�y^/l`���B�C�|(���>H��\3��\
2���=�M4$��A�*9V7�I��ޢ�_��d2����O�A��۳�ǝ�OlO�D��Ʈ��5�=��f�u'�.��x�֎�;.F}�u����k�����A�`w��x b3�I_�ёC��<�1��a`nmm�:/
��U�� �%p��~	�nfQM!�Xh~���t�4�̟���t$] J*��e<(N���H=��X�S�e{��Æ��([�7�1փ�V6�]�}�?�R9m�2,y�9-X:��T�����Nc�K�MM�jY2ɧ�罏����a
��a���^_�O��f�stt{J��f4C��}�c���0I�I��ϊײǸToe�����)�'gU��#n�������0.�2�7typ�P5j�Ǩ��]nP�5����0�(�[�!�"���Y��K��0�6_��ɹQGI+���pRIO���
dG��dC\zM̺���>3��r��N�Ȯ����+^� Y��|��b�@�z;H��L�4Z��eɲDZꗅ^����$9�C�����g���A�"k�Ns�ѿ��$���խ��<6cEl�@I��ο�_�h��c���QQQ������^^ԯ6\�uT̙lll�Ν�+�-f�tQW�nR������Do\%��>_w�'�%]=��ݸ�?mI%o�����4��"5��n{!h
��cH���N�f�d �HՓ��u�^u�п�=�|(;ZG�~Џ�|h������`�	A���vI�%PA�
�CAA�T�bR���bEV����RM����K\FFF!���f�؋KK~Ж�H�#ŉ��QМv���՝-rц[j�R��$t�a���{�ܴv9�9�������������M;�Y�K^=K�dN�H��EѪ��	ǻI��}�v:7W�<08h���PG���B]I:6��x#}33�� �?u���f�`ӎ���t�T��	H��v>�mNΘ��mN�nAێs��_�Kݮ�1���:m�8�R�i0���+�z��b<>ϫ�r��WK�oE;���ܖ����\�����3�_B���l�%��e��2�`/)���r����=��0Z�P��� �;���#+z+*��<��rvv��I�*I�%<#=-8�#�����mޗ��kٺ�z5�7�h���skk+N�r�����fw�͏V�~��@O`�:�����|{�[�n�yT�P��ʓ��e��d�q�4�Q��G�嘰3����E���c�cs�D��
Y���'������������E"	$~~~/�J�D��0Q�����ݤ}XVV�ߨ��Nx˧�c߾^lp2l��F�����t~[	��Z����zǣ$�������&,���տu>�g�*3.�b���cr/���,�W������9�:㸃�Ŝ�tF�~=Z��+�
��!�<��S�Ў�U�Hq�;���J�ӈ�h��m�}�R?ve�~c��j�L����ӭ�T�}_�y�3qmƶݞ�ؑ���]�y�Ƽ�L��\)��ݱ�77�F(^����eV�egا������Z���sc��Ј��0���`U2�]�,��<,.�x�������b�	 .Ao51���mqw{�*Ŗ�PB߳�K��SŎ�
��B��h��}UT�W���@����vb �ut���O@������������u>�{&���R�ې>��}\�T�%t��	�ɿq�#�/�̠Bl�E�������u���g�L:i�7,���~+�p#��hv���ߚɒ�C����d'�֔�r�#J��\��!���ɕ�իW&����:`��L�������z�����mq���3���j�K:f@�Z��lߦ��U��.���z@��w�؟BM���G�g��_��'Z�)�{|��'��Z���3�!R8���-H��s5���[�g�P��b�cys�nqO�KZx�ǋgg�m"a�S�[ή��Ӌ�X)���^���NT��v�S�6&dXk������
�W��C4���;v�	��ʽF����ND�����EW[[�_�z����H��_�pk��[L�b�/�L._�|�ڂ�:1��`7m�K���,~���h��o���$��#Ƽ�?=�,��lV� ��v���y삢��z�x�cN���iy2�޹W�O&���5��%B��Uf懆������s�+�x:���>���O�ts0*o��:�*���w���WSVl�$_��Z���׿�s��-��8#���Vɰ��y����q��8y��+󾵶����u�������6W�A��$�@d0�v+�cYb\��� }}JTO�+(��Zi�:��	�AC��H���r�W�U��6T��HȾ��5ch��^����)���
Z6f��+����:_4���}At�M4Jpsc�s�~ ��߾������V�i�/�����D��=��R�Хy��&3��ߧ�����OX�d�o��/4��� �Мtqwg�,Χ�j��[���)/�i2O�eI]��~��>:����bQ�=Gv�`I�~+��uj�6&2���?�1�=�ZX�3q[��}h��Q%�c쐕�y���Ą��U��4��*�#���>D$����.<e��F~�(.�ڰNZ�d	<����$��!Io����7��ɰ��d�`ɂT)�v?��{܎�(0��j��i���N�e8��H�%1sHݟ�
gz�w?)����q+���$�YTGPo8�P����#����/XYgC�0BzkCx�n��[�_�yN]�V����MS;M(3DTp���f�^i��Q?WT�c�9C�m�"��$;śӖT«�ot�z��ڥ�h��<z8���\⛴�!`5�Τ~ݦa>_�=�]��>`��cG<ݟ:��Y��l���r԰v��a��i�	[;��������46�'	�W��J4.��� J� ����������-����S:��V�5��9z��sD�-��qF�/p��
ҫ:we҄
� ��י�ǻCӹ�� ��Fς��0�m�3�Ѹ���ˍ�����I���h0�7���V�iӣ��>� V�,0h�ؐ�u��TT]��̵�'�wH�O�
�/(�������{d��r2�wT6��`�@���-��ϣ���'�gꃇ�m���:�l�f�L�fQN���}��}���6��� �����g/�7:�E�n5��b|IN~E��?æ̚����>���u+o��$�E6nr�TQP��֚��9v���--�9�/B�_����>ο��9f(�IHI�\\]��X?*�?ڢ|��D��D��֤ۀ�%?��&@�n�����
�.?��A$
��>&����Pz�F{yh�n-�S�4���X�Ҿ��]$��1�&����֫Jr��mk���Ƨa��οv�1�~��3��x�E�W^�=�Ha�����T�P���H��%���1�������m݃�wl	�DÃc�cG7#9^L�˰��o.0ԥQ��(��v���\��.��|od�,�h����wO��dL͋�|+Q�ѱ��E����w}����J�P���Q?��"��ƺ�}(ℎ���N��ܺ��;��͗�(��֐��ۅ�s�Z¯;\%g�M�)�oξ>��d�|_A���(��;����z��5T�� ���-�?B�D

�\uC���D�张=ApJ��g�]y�Rgf��H^C)���9A���o�M��X��~�e�~������>�.��EDZ�g`���|�G�=�w��#��vA��P���S籫������c�P�"��7�r뛚�FS��}/&��>�����iOzzy�.�e`'��	���+���Ǽ�t��:�3<^l��`}&��[W/��9u���k����dP�Г�*���g��N�X�u�?(�k��\��8&��V���I�;'O9ޭ���)�偂O��/��DFJ�L�(&����N})J����|������ ��1�9���x��p����++�3�K�_�y�r�4�R��nR�>(5S�E�mE��� �ӏ�`O/�ө�]��<Eq
3�H���%��؜��ϐgx�I�e���Ͳs:3E\s&�4lmn�BE���>Z?	@�8f��/����j���Eg7�v�~��]�Z�6������)������8s��}bq&���}���%q�]r���`(��q��ܪ��+)--�#
���Ύ�Iv66:�&�V��$�`[��[^"��\<��m�����@G�����$�o��s�=dcRF�j6�{�ԉ�h����7����Z[��nܤ;QSF������H�pTVV^�bn��X�2󶗻�9;7G���`N��P����+���vM�	s���w="�7�j��y�z;=
w�B�s�Y�J[C�_�d���د����O?�YM�0�#������ݺ2,�⛉�E��z���r�y�����M�t�� ��~���dݫN���o.��؊R�����F��K�����P�2=��s����涻�(֖��X��gj|k>.c������,�	_]`qI�H�&�U'�ѣ{7���J-3-��4@�]�R��5�������i������/��=[ ��<[����7�?ZH[���]tv��O�B2v�Bؓ蓓|\N�ܞ1Sct�w��y�m����yx�
ꛉB*�/Z�$���$�w?|B�jGr�r�X�����)+s���N�XA�Fv��̽H;�"$ ��GEe+r�{s]�ꥮ%{r���Q4t�������؎JD��+�v`;��J�A�l��(����1�[�ﭺ�!�,����+��5O&|B޿�HP���x0M;jc-�fA��rnB��hB@S��'lՔ[�	��J��"����MFg�\���+q��w��f����]�a���� ӌZ�ɱ�x$?����wp��m .���]۫��2<q��Sܲ��3J�N�m���j��ލ���bh/3^ޛ7���]+�����M-O��'��,뿖=-�������&�����Ǉͫ��Kb��l��eB���%����\�ov��^�=�#�`G��|l}A��t!9)�?��EV�KX^����Y9
C����u�f��-����߷�u��N�����&_f�%���u��5Ty�9�nU���#����K.�Z�[ŕ����J�@���e��4�����d�8f��]�3�@5�qM�<����Į"���*,��.�^b�#j��Ee���Z�������DMEI�c=Ĳq,��v�)��kE��?�;hŴ����浽�|��{��y<M���(���X�vH�i��:Y�K�VV��W%�ex%s�?�l���t}:���8�uIe��L�O���'��(v�A�[z
�dt�xoм�k��ۋd,1[�����ŧ�|,~�#�Hs�s�<S/���|%�gE��b����>ө|�G�/�,T�Q�dO�O�.Hk�%.�7Y������]hU��Y��gFZG*� ��O6h?�^�`y9re` ��0"��v�C.w�mo?Vr�vH|B�M?}6�3/��mR\�m����#
��f�ya(��7(���T��Xr���d�q���t���NR<�ƾ��V���?,��� {x��)�����mV��F�c]]���y�99.���{�K3S�z�
ߒ�hF��_���;8|+-��0�C�x���2���`�7R�[�(+.��
���o=�0���������&:��������qc5H���Z33�nί�鍱�|��4�q�c���>%�2t������`�/!���k_��G��F:��1��(�j� �z����s�ej� ��������oՊ�'���tZ�91&����ܭ�K�Ӿ�����͖���t������:O��x񼰶�1K"�`s)ij�ċR��]\P�1I	$zVZf���ߝx����Ş��,��9��1n�R$S�)��urq��7���_k5O���A�ku�����Ƣ�np�m��n��t��晈b�ݷ9��^�����F�1�eO�ץ��jU(xL�[�sp�!����`������*.�$��5呫�� }Ɏ�������=��ʮ#���"��Ks��6n�����dV�vz�}�3�`"�(aS��������$��"�ق�fzb��}!B��(+��/�3�ֶ6���J��~���r�O3?/�A�Д9��P���������_��0;N���ԁ�R�����=O��%����v�fh��z�g�����Eޑ��M	��z� �X�re�XyW峛h�%])�����q2������~ pB�a�����\���(q�����f��kթ/�j�==���!Ls���Ƅ>����.dX�v��l5V +99��JUV]Ww`L�F���'������fMp1�H񒧧�mj�h�`~�>5u�[:pG����Tz�1�W�2�+�.�ۃ��l���*�â"�Ҝ~3mm��-E�돭aE;��M�H�R�u,��0������3�b��95��_��A�xq&���?�J�4ߓ�R��9�W�k�sIe�7S1�:�*�Zx�H:�#9p^:P7����5>�G������K�\e�b��䯗a�8�j}���9j���Gc�`��ä��t*9ʭw++P�\�<r��[9�9��C�lI�_�6`�dgD��f��t	n�������Εv�zp?0}������h��@�@�ԕ�K�AG��g⧻��P�s�������]�G�������&�ˬ/�>ٙwEu�b��L�f.T�A�׋�F%��G~�&�zF ��m�/y�����߆=~�>�~DD�^4�.ߺ�����bI���6��盬q,�W�+ZKˍZy�X�&����:���������l�x�k�&IL�57_7}�D	�H���ã��t��ͅb^��}'����40�}4]��3�nM񿦲g�FxO�w�0�m�~�#��?>o��7�;�?��UX.�Y��B/,셍�J+.��^(A9	:�?�ts2�3�ބz�
7�A	D�&QY{�$[�%��}�0�-)K>�]�E�X^�NJ�%cM<r�5G[� =�"K���ө���(����H���\�{|�O����ii�74� �m���sz��r���Z/L_g�)x�~���$?�ck��C�|.䲓��wP��n7o���f��Qԯg��C���!���T���,;j{@ ݯ���A�vr�� ����tݎ��/%�m�b�����x�D׌�,�C�ǜ�8�le�-VWs�<����0����ݣ B�P9T+]����f��i�c=��I.՝V\���6���(���I%�P�l6�:\3��������C*MۮH���b��'���&��c��|�e�{;�s2����NO�q�L��!(1�ʉL����:8�/c����C����jn\}�J�}�=���_YO��O�vWG{T���U� ���c%B?������$���������vH��9����7|!D�����6#[�<���#փ���Ҩ��}in�7�?<VX�^&V�p�|$q6FG�`�\�)�۪MU��Tf����JHHL��Y��w���On?.�S�+޶�>sn��a�G�7��fv����߫߉���ק�7<�%��E%(��D�]
���nl!Pc��Ò��£��4�J���:���2�h\���3Bj�����_ۊc�ɞ���+��N�L���r�����[����zD+�>�9��?��8���$544|DI&k��~sqw�Ӽ���Ǽ=f�vM����X���p��LO�~����T��������_�Hp/��b��Y$)�:%�i��P�\�kQ]
�@yu7>�&;��7�Y?�V�����Se��q5��JGT���TM��)�&��@�b6Qhkc���#Ո�(R�d���i�F��N8������o���$��[�5���,,�L ����]v�͈���`-f�)BN�<m�ۢə;<ΛT�W[�-���	['P����Ėۏ�|���I�2�����7�!�q���2CS	>/����u���?`����E4|]_� e�=ɞ#C��On�������ٮk����/�Z$��n#�lW�d��A��6�ژʼ�9�rX>'��J�+e�k�׿���o ��!r�x��/�o�ك����y'}���|����ɩ:,�We6Z^Ց�b6��C�ch(��`�D[_)�����s355���!m�ho��Wo��0^�c����ʸ~:1.��<���5��Yv��2�f���A����c��f�{�7��5� ���i���8 K�/�/�ftU��ᔼ�3������y�ñ�s}25	j�E�&"n���ۛ7��R�����h�B���>"}52N�����t���jU�qS� :��e�Q���"��9�������`o(kg�$
*�6�;F�ӕ�C&~a��C����^nw�^̝@����ۜ9��F^��y�C��W�E�]��T	N�$u���؃�:k��5�4�����H���䟢���*HT��F13��0��_�2`JL�ڼ�� ���fVԛ�L�Ͳ�:N<��.�i�_q�b��	�]�rz��4;���K����uA������r�:�5�x
H��j�M|�����Rt�$7�@~����Ģ��o̵����<A�=��Y~Cy��a�<�bAnp���*)�6���2ǖ��#�"����ψ�kkk����bm����o>0sW�װ�=��"r?ȀA�W���82ē���=>��S�󸪫K�\��i�_� �N��3��߂GTx���g�������a,�r���U���P�N�9-�Į�>��6���Ά� �N�0��B��sh���;�7���6Ø*��a��%f˿�Ԧp[!�*f?�`������L{��P�\Y���_�����˷���*}�B�Ho�Kv�@�ƊԊ����¬,#[��oo���G�,��w�K�Y����z��m2��W��},}ss����S��5��2r�����%�
�(WUԤ�6��I�ڃ�+�����W��36�9���4�2�����@��F��WL�vۗ+�)�:��59���o+�俗�~]E�ڻ�<�a�����J���>*~H�q u{-*��l�;�}��U��M�"Cr�����������Ne;;�]���Ӯ ���?1^2�I���{G�;�O-���k��Sl��e�W穳;��������)��Ε�
�W֤���T�u�X#�Y�o��b�\�/b���q�ٚ��hD|�ђ��%�sW�k�|6���5ьUŴ|�uAr����5��/��W�.`�h����ײ{xPz��Q��xA��L�p7�����hmuu(�)�%�&|5�I�ĘP��JΜ�5w��iwyl�F��edP�m��)G�j��ٹ���-�*�Q��TP���z��8V$iQS���2a|��Qr���%���n�s�9s���Տ��8)bPg��7/����|�"��g9gvE��b3��gje����p�-��|���+72����
��6Ii���4��[J�#���%�^yzUq�6�(�����n�:�HR�.!j����Q�ԬW����pFEI�����V*���?��S�v�|A$�/�������ls�����EQ��of,]s6�ak{�r>�R��X��m�!@�l�����>}�4/���L��
�p��ax�/���P��:'����p5���hpd�Cʝ��"p�q��A���m	�B���ƅ�������T��͏H�()S�=Q<����TC�wQxd;�����_�?[��<��@	=�Т�\��(�� ��w������Ʌ-��C&���$��t$�iX�,KNxL.�LJ���1�߭w_T�@K����"YeE3Z(J8��=��cw[�pw���T�7\�{�෿m�$?��.�ԶM�`_&!C��m.7*���X�t�84���9�4� �sG�K�)t�OâV-
�5��"_���a�-��thE�#[I~1���_���<=~H���L��Ru"��^`s{���y�|���9�U�e@�v6�|Rt�n�J6?��i��ܨ�b
���ɮ���@�ަ'J8s%bM�R�RP��ç�=Z�$si��}��#���[[[�֧��E�Fg`�A� ���O���)ĨLB�<��~�@���B7���d0���7�UJ"��%�}1�c��q���T�T��b�� �y3.��y�,Ϭx�4�VU#B�`;��ձ��般�
���P�[�xL����(�"(L�o)L@q{K i)�zI�6��jO9{�J�F+�������)��9� Oϱ�ǣH7�f'^���OS��$-��v���ٖo->MH"̚�V~���#�<�ʲ�r��p��`�ό�\�.�Ǟ��^Z�JI��r[�>�E,�Sbii���oh�A���tƱE�M�x�gvuM$6]��?+�'A��~~7L�а��;8����Q�Y�N/����t�mP|�	8ތ	uF��d!��-O|�� �3�ܧ��_��?Z�������d;�Y�ƪӗf��T�u��+�m�6-U��c��QK�q>�`�z6���i��?�E{~�P{�_����y���{ @Qq�#��gIWC�2Җf�.���"*t��p�i.%%�+�����kgeCC)��С��+�^fn���5��-b�QPtw�yS�`��-�B"�[)%�%e9fj�-�5s�F������R�1��_/c*�>'��\R	��l�Wf~� yڿY�v���i�ٱ�p���W��9�$8�P�֚��4�u�gf5�\���ư���ҭ9�e�Afr���ݟ��2�G�|L��]^�*{A33:S��O����C���]@~��������.�l��լ����;#���EKK�^�ء�YEܜ�y���$�_���b%ă��%�_}yL63��x�:n"�2�����=+�^�J��-�@M�x�Zn9UI���J�q��kSX���jl��y@��&�q�4*����_8�~���=�����5$  @y1ɀi�����?;!--���sr\P�{q@����x�n&���y�	k���c�⪣��70ϳi��n�B{���G
�To{��_�ok63�*7@�/�'Mۼ����l�SN�I��z��03L(�����Sx�ے�"{�f�hW��!�{-�� ?��;/�18���D������֟���R��r��P+����_$.���s�ׇC�GI��e�1��~V��L~W��09^6������B�WT:�f��'w��?�R�2�k*w ;�~G� ��^��Uu��U��b��*e��at�:M[� ����X�y���0t�<��ho��JJ���ֱ8�gJ�jp�J
	�b39��3����2�p]5�{m@̧�ȗU���|�!��Z��Z���̿���~�CIȢi����FOh��D��=_V�b@�mkm�q@� �e[i�xXǬ����S*g�^�շ���s�Mb���IͿ1��Þ���gZ����}���4�\�~w�^3*=�ጜ�ܑ�|��X}Bc�aل����.�� �u�5��}$(��O&%㽿5u���4~�z�})�?��.'�aӓ���[	Q�茘S���1{O����-^[���c�l�l����E��U��f�&TBI�2���n)],�30pj���&�wN�!�����_�^��o��W&��8*�GLO�ª��CL�m�͛�~(���U^yop)u�)�{�ڈk�k�̪NV�q�}����LK"���T����ד������ll�c�H戥W���Dv'FO��bj*��.J�Pt��rD������Y^����s�y��C+�Tm���[�A����e>�%g�:��9=��IC�~|z�URJ#I���j�p`���3�L���*[��ÌE��W�Zf���0t{�e4��ZϽ&.{D�/bZ�d�p��K7���d��'���!Cୱ���0�������j�<�����&Z�����D��_���C�ℇT8��0�.��R�s�+�Oqvv�n��2�.�f+Qs���a��\f��:E3�I:	���$}�^:������Ľ$�Ak��X���ό�+G�SR�u�ט��~�[y��ܧ�6�,1W�ޙ��u�U�e��ßWj���3�Wh�,5�۰�6.��]KO,*	��l�'b�*�T��l�I�R��H�,��C��=/��ôx�	_�]�\�`r����( [CN��6q��H�_�C�މ���P�(*V��ױD��C(2,Aw���+�͉�;L�wNCa+8�8��?���v|�1_`l`<&��ϊ�NN�|������N�ƻS�3���x?�ջ�>&[A�){��y��R[@���lŜ�~r\r�o�\j���d�u �?���k.��$�~�݇��,�WVV�������|%	p���:+;*__zź��*��<|�o�����]LC��T���u�1��Q
T3�! ^�~����tSǌ�$jvbB���mtG�tCSSj�g��VUV��o�^�K��¦F��V9�M8�<E�#��lN++��f������*^O� z_����*�i�P��~B� 
���um�����&&�pY vc9s�B ?����M_�#�yn��EKBwpK%���]�k���g$7�QL�RUR2��������K�%�ebȧ;tߧ!�@H�Mz^U��B�Q^ۦ�m�X�'`Ҋ8���J]�2�T;Ӽ�-/�[�u�W�G���║�:S��ӭ3I��0n��lߩ�� ��C3J�c�Xf��~�1;���Y,.?�Tݟ�Jm��'����ou:@��9�R�*��=�Ҫ�&���zi_�b���}߬��Ĉ���k�]| ����P0���I\���/ �CZ�`s�O}1�B��G��s�Lْg��T]�"RL�=D�|*���1��uu���������p�,q�4���|*WR�íM��ytI�z���JP�U�~�L0.�2j1k�jg�*���/�,��VķX�+�q�t{;�4z��W5_�+>�R�+YT)��PR�`Q�)z ��Ly��/ށ�Ӳ��?���O�د�h��H�m��츺m((z�b���)ȳW ��4t[��].J�����R��ԍ��������풤W���b,���v6�P��u���X-'~���A�w�O;��O:�$�X ��	������B�?E滕�Ԕ������JꏔǇH���Տlo ��A�T��sF� �g��F�0� �rfΩ��A���s��B��&ب�]E���G'�0Lq�����Cm'U˨�����S�bI緲!#�7olǩ�<O&��@B�z�o�~�q�T�.x[����YVY�k�Jw�� ,
��.�p|g?�ĩV}�++5�r�=��c��e�/�V�5�{ 7|G6qZ=���-��m�<}a$֕��Bu�̗`�!`��j�(�#e[��t�To�o�*�%T��p~�Tv���eD��NU�E��� V�yj=���=�֎�O1�>`e�����������A�VV4���Yo����m+���ȴy���&V���^~E���7��Uݡee��(�l=���e��2QR�ɪ����b���vW�p0�l�F�J�����ٿ$fd&� 8�F`�ޒ�Q���Y�{�L�`���F�%�ez�o�LM�f�f�GxXD����=�%NT|Q������(���m�;h0��s��¸2e�����3���)��X�tТ�j³��@�cy��ȥä�q��� �����4u����zo_5jY �
k�.,U��s��_�c����[�<-��xCɣ�<ڃo6;u�|�kjZ��T�ho�UyX���ڦ�}x�[_���e,��F�\x���˳�()q*:.ۣg��y%��C�tA�޻/�������jB��5.?��_n�U�zK�[Y�͈Z䝮�.�y>�s9�/�Ue��yu�w���Vݳ��
�t�%����"�08ȑ���.���/�1�+S�S�������<spmWq<�B!���������ɚ�Z+��f���p�t�&�
-++C��Sx���A�2�
W�W��f���}+��9❇�IQ'*RΔ���2�{-5\[�.?�n��m}?�}���@�uFLf����g�T���;m�^F���U�>��~�f�Q��w������xfnG#���|蹝���W_��^�Np�������Шv����ݕۑ�F�]�y�K a�p��`���<s�пL.�4�e\�Zi�v����6tpp�� 79/	�y�0m.x�[Y�4�>]|�<R����B�_^,� S�9z��ʕ� ]��T�����W�ZVC��K*x����l__��8���6#�P��An>(-�u7oU6����8�=N�����	������6����QӼ�dl�pe��Ѝ,���� x�!����gz�$R�:h��ِɴ��ͅ1�d�*Q&�,K�	�svW���iy��4�n8���@'\��e�2}���s����1���U�<[�	p
������_n���rA���A�pf��ۭP�66�B����,���9c�֫W}i\�χ�S ����|��v�}R(<�\��O�� )`t��� ܵڌ�$��6B�]��TɄ�!76B[=�����_a�p!f��*�Q2"�h�F��.�߿��POW_?^|��|�C��V���f�yG��S�dI���7� �w�N3׀�����?���(�����X�X~�K+@:�uF���eؘ�`��=��!���֭��RJ
�
�ՔSq�&[�����G
X���Z�S*W�d(.�;���M��1��+�.�h^��ßN�5��p=x7�� ��%}j1..N��Z�e�e7��
9�D�?%m.��`yͷ+�Sw�[x��#!�yﾦ�I�y9��aj�DW�7]�n����X����O�->l���� �۫]�[�S�c/�~�jM�\;9��='V�Q걯�b�b`d�}�X�,Q`\���������ԨN0(�R�΃����/����8��b��s���|Q�{��a�K�������	�I�%K�d��n��A�ɾ���De�NB�d�3�����u0�d7��'���������uu]�����|���r���G��oϣ{-��ycN�ʃ�����'� �IW2Njk��KB�e��ئ'j�f�X�D6 ղ��DD}�<v��!Z�2#��wg;p��!��Qi:BTl�����;k�|Ș�ʊ��W!`���c"��.������k=�������a��7Z�=Z���B��m4��&۩�����{T��S�xM7>�8Yb�;���'���%l�J���G��������Eۺ��F�3�f�;�?�%����e�1ڟ!�gN�81�
i1�I;~K����+ל�����i&l��Uu����
�F�9$�93Ǡ#��Q�K�I��݂��L���������MWў�G��rN�e����h�M�H��6�(^+^�*N]����/G�zꗣE�׃f��L��2~�)!�b�&"o�Uydqqqa2�\�gr�{��!+�dp!��J�v`� ��Xi(�4�Կ�{ez���Q��1��5E ��Ѓ�	o����5�|ʵ9r-6�ߟ�N������#f�W����,U���so������*�������)��U0
�~u����C
v������F�0b�2�6)U��Hc��#��]3�2<�|4���;��OԜ4ߜm"��ý�+zB���\����1������?�;��s�k��N4e�t��}���=C��V��<�"P������s�W����N�M�Z!07��\�\����tbg�r���UCi��Qd��n|�֭�|~�����WuƇo�@�YAAe4-��˨��$����b���1�\��R���Ma�'k�b��\swM��,%�t^5;"�C�*�W�J�&0�[���$���N�KH�4����/�{u�W���k��T]�*8u�ՅEw����C�Z�h¼Sr�����?~;�Տ�V����5\��H7���4��f@�<��ܡ�5��`�f�Ĥ����/�[SRa��2<��K�D!A9 ��jy������w/�´Ȳ�;��.c�fԇ��ۃ��`���a��h�v�3憴s86>fQn�*���r�sqX�U�(+��u4�ݓ��A�D�2&���/
��S��M*��oaQ��^����{�_����3T�-O��$I+�΁�@�8Xӝ �(��eU��kcն>�.=���<:q����ɳb!(İ���RZ���@u���Md*S,�6�dϳ��f��eọ�SsX}��q���'>6x9�mS�I��)(L�*1%��d߈���Yݬp�:H��F�R�1�O���Á�3�C�^1�
�v�og��L�'��x�~-U� n:����!&��ƀm�d���K��)� ��Ҭ���<���3gΐ%a<=}���M�H��������:�<�)��妬e��|�$'+^�4������䝞V.�$5�Iv�H&��uf�#s �cU`�/nZi^_jb%��e�{�O����b~��,�
Z����\}���=������۶�dIsՕ�EE���U޾ިQ�Q������5������]�c����{3���?O6��A��Z뺳>��k��ٳ��� �Ib�ɟ�t����ݍ���vW�V7ߴB�|��>h}��<������<��Cg��Q�k�tY�����`jw{5h{���������p���Ot�Ehߞ�
-DA��%�=��/ �����cƾ9�B��L���\�Z �Y �������-�%x1�>J&�p�`.|�����2#f�I]�c�1l�/�o��P��q|�������ִ
�����'F`�b�uV�ɂme�P&��ً|�/xö�2��\��|��'�#d{{�8�"�ţ2)��x�Ǐ��nSC7n�x����=<fa �sX<h�v��T��[~@츬���WVT�d��������|4��@1��]/	�v9U�8M?�Ʃ�������xv�i�����z��'���V�ֻ�	U8^>�{�m1��|&���?��s���^�,���ZT�I]R�ϗ6ե�5S�~#PNAL�U}{)�)��}��b�*�i��2�_H�{�D���J�+?��]h�Y����0*aLR����tssK@�c��E-pR��C;�ڸ�v6F����Iʹi'�wem�d�B�A)���V���Y�% ��HB���V3Ƚ�1�4��n�߀m~�o_�ᒲmT��-4���;�]Ȗ���o/Oݪ�4
�7��>Īr>k���W�o���O���"�S�d�4��څ;ߦ-Q��Z�[Q7������U�P�G�viA=�F$o}������Q]�j۠���^�Gӟ�d�ua�^�uk�>kZ��j&�;Q�K�cI���۱̡�iH�����p�d��M��^íJ���z]]ݭ"��%|4����c���T����Р��i��RW�r�}�_Շ�Z�{�r~Sw�0L�@��D������DDp��y����e�6�^����I���Q�JbCl���ö�º�z�+*+�v~I���(�%%%,���$�Ǯ��}�_#>�6�)�V�:6������B�}�~}�lonR���|��c'��D}c�$��z�M|;�yA��F�h�JƗK
Y��Sg�ڻV�c�7=���V��C���<z$;�z���>@��������߱��=ǫ]G7;a�i��q����|O��Լ��ժ�^S��ND���܉��sT[=klb�Dy)��c�j!a�����}�,�ɫ��d���m�5�����k�S�J͊�m�z{g���qGm���϶�����F������N��6�Cfo�u$���������_u�8�R����/Ϧ$]z���i�Bɓ
g�ڨj(6��5\����X�+	5���K�������ߒ���m��_sf�.��<k�3e]�1�VG�#'����d�V՜��EW��B��ݍ�"!8��R���q!Qq�-,6L�b��!�Ce�{���&M�W�I{�r���a3b��W�(?����������Mq�'���3��T���á뛄fah<��5V����(��b��O�p�bkH���_����~Lw���җ�]z�F��s% ݦ$�M��콰��;*�V������T�%�e@H��3\��]/��h��҅�%������V��̓���\S��[��k��Sh��y�A�k��e�JX�~7�H6��� �����V�҇�iCC�p3>�m��Z�lu�9m��J&Ut�-(��M��7j��P�d��*��L^�`�8�������R�BW��ȵ��1w��G���D_ԑ���3��^��3AAD�w�USs���p�b��� x�j|�Ph����*���C��...�[����I;4"�l��  �*�gm����%��;3��>kT�����(�Q�O\�߾��+G�+�T��[9ef;;���*v2B*�Z�PX9� �[M����V��jn358b����,@���a�p#��䧡�~f���? ���Mc�s�WcV	���:w�vnݓ�9j$Z)���?6��5 �D��ԩV������� �z�/��[;�̥���ߊ(.^<�V��m �����r�'ʽ�f?
a�
4�����zP���p��ٚ'�����V������YA�'���.ʷ�b��MT�c�O�}������em�r�a��������Mp���Aa��A%���� bq�t��G ORs�$���w���C�j�Sa���$&U	�}�0���̒ [|���DO�|���������tp�c�Z�O}��;��C]�an���y�B���pG4�޲j�:��E#j�OR�3�Ƈz�@�Mv�?�6>l��h��`����I��ĩ�|�&��i��������XG�c��b�X@}��d�B�7����ۣ�)���̋�c�G� ۱@��`��1	<|��|��#<�>p^���ą�x�5c��~|���L\�!vc�5ڍ0�	'm��ߺ�\�f2�l!7�Rj��M�+'''M���7�m�L��� ���>id1��A�~��x5�ݕ��5��i�(�ٟj�f ���L��Q����W�x�S���1�<�}6��xx:����b�r�㤿�ZIn�-99�\	v0����Luq�J��U,v���-0ͽx'��9G=���<Xs��DA!�,J+h���T� ��76Jڽӧ�L��� �o6��C���|�!�HB!��Z"����db�~P�R�n�ݕNp���[4�$��'��Ò8����� �%�<�mwJ�90p��bc��;mycW�|0�d��/�,�!"���q�;	I�cs:�k�4�\�OT�	-v�9C��4M���]l���FH&�m����"� 8sQ����w>�b����1|����dK\�I�Y"�8i�~�!�V�����0�C.~_t�ݺ����w[�kR�	���]�a�R<�A)���f;3�Q�W0vY�JhG�%�/7Ū`&+��f`������%@�X���� �H?A��bQ�)3��n���|�YuC�^�d�w����)�UW�b��'�Z���b}ұ <?�TM?F��m���3��@��̳���qx��h�hW��vk������������(Ƭ�������lu�9���8n~�J?��EDIY$wT�s���lmNҒP��&\��8eVUT��"��VV��	j��������y�^�v�p����]�	^��:�D��?��q�Êq~�ԭ'O�<�����EN�`0�	 ���4y��0:�H�=��s��Z|�q��8YZ�Fj;�fjb�W��jfR��upJ���F��׳!%/�C�o���{�V�M�����7W��؎]�1�������%����b�)�����̡��V�f���7���H�`���=(o,�߉g��Z T8���\6�l��;9�&�|���wv_u9�i8i0�������8 5?�4�^��«�?��1$x&�Nj u���M�q�
�`�,�DCc�F��b�a��J��s;�4݈`R?=IWW&EfDv$��e�Y�LĪ#�|a���9��-�ц�	E-�#a3��M%a4�P����:A��Z���%�c�|:���&.A�Q�vvq1:���D���� ��+�x�\�1���-v��t����UI�@��&W�G��h
 pQ0��
�dV'�D*�sİ�(� �h~����	�_���\��_T�]�'�~yz���R�i��k r���SA�h	3�����㞊�h՞f�S+ܣ}P+'5�E?b?(��pr�)_���A]�<(�\����S��0���Q�T���2�}1-�!�=����mQ�p����-cSh��G�y{�fM���^���,��3_�E{4j����"��}��B�ٚ�S����~��J��6�~-Wj��{N.x>?o��P�t)�����Q��;&*YB��y��w�V��
{���Y�a��Gu�%��6��*k<N���I0NU�J�L��[,vbPcK[�nmac� �P�01��a���
�\Ex^�j�I1�(�?�{%���"�>������u�g���O�^'�u���*Td��n��v54�a9����ݽ�5IL07,8C�XA��%�_��{��~���_�	4�;�������8(4�lg��7���Qw�M����S�˿��^���i7$�k���l
k �o�mHlj&�T���@�����j
?���� ���&Y�b� 	A�ݒ+W�:��� �N�����8{���Ι}	�R�;s�V���Ǐ��/�Y�ބ'����>��8�U����m����ml�0޵*;{<6O/��Ԯ�����P�X��I���Ͳ�Aot=+kՌ��;q�e�5I)hͩ�|��]�);���{{����Wtڿ%^0���W֚��SNAa���ýޣ�\����:�.��_��m��O[XXT�%_��GH	@6;<�ι��ö���<�~~��D�V�đb�e9C�ƞF�"o���Y����[�p����8�*l����7`�T�}�'��gj�������C� T
9,LTAo9~��~�<<<������n�����͇�1@.���^\��F�,��:=��9�V>Z&.aY�������o)��gX7��`t��MyH�ϟ?k�v�g�d�Ub�?nt��[�*8G-z���A;���� �WE�s�j�I�*��m�c�r�S������|�WV].�h�&)��P��1p�ǝ���Ұ=���#$%���45�_!ZEI��DeS�hRkg4!��׍ot$�����ڿ�e�ȣ�;[�I�ځ2���F��L9�[�0�UUU7�W���Vi�!t����S(ҧ0��R��Ӆ�g�@�+�f �B��$Hͪ����͸�%�����MKȇR����O�!%�FJ�GZo�G~��'l{���K{��+�e���]���[N�Hr�t����bg�`�t�y>-=X���v* �a7F6�{7zkk��;rz���\Vv��j�z\�m^bj��M���쏇�GL�CH�Ơc�^���x� �n�J���\{�,����蛠��Wu�.���M���'n����Ȅ�_������J>�X4D�3\�p=�5�����g��C�U�3�I9j:�K�R$Ҥ��Ѱ(�����5W��8�ċ��QT�_0�z�`���cftw�R�-�`�OӸ|�X�b�f�HWh��
����_O(N�I.�ͤau(��A�`w�S��( �?G.!����""B�!S��a�;� ݀����c�[P�#

���Xo��G D���2�_W����J�A�{�}J���v!M�a��aP���{��yG��/"��W�����~kl(�2��K&�����pY�e��]ɻrE%%RǏ�����.o����t��kE�E[�7d��72b�;7??���_vnn�����@nOPa�-�+�\,����T��l�$��R�&����u�Ҳ~{JJϕ�J6�����+0�J2]��`�����r�66�Syy��"�`���V�`�5�(�!�.��ٞ���}�F}t�P$c�-e��R��X�0~��j�!�������?z�ԁ�>M����_��~%P��p�V�z`�n|����ӣ�=�B��AU:ڛ��?�N2ls�aV;���t�#����io���
2����@{.�5M�Zh@Md��b[�	0����$�cX[���s~ºo�e�$8w���s�/��f(�ܻ��f�(5���5.CM���P���3�raȫ��.ϪC=�{�#C�Zj4��VI=Nhх*+)YA�ҵ� &���	TE�싍p
E��N�� �q���ՙs�Ln�dG�?���\RNr2;�b�3�Q@��U3��;�~���	ϕ/�~��o����yX�_B�8����O?.�-V�G9#� DX��PuT�\��OͿ��hZoh�;eww��x��N<���t�L|\W
���g:tC�u֚o'f_�FK%�ⲭŤa���f�R6�F�0S���r,$ڔ$�[tU�\[]@J �<H���|�'3��nKZm;>#&&	��(�4(8�#²��߮��.�K��b[�,��,L*_�R&�e:���i�p&�֡�����@/����q[G7̒�nv��!������IB�oH���p&�6�Z���O	�+((�j"�ЅM'��q�J�:rB���GI{Da'
�h���1�
�w�V�b�y�S����>���N�e���s�����Kr*bX�y�W���O�cd:��ۼHL�q�L��#'K�Jꐁ6ևPE�k�o��֟5���@o�s���}�P�}��j�LweN&cا���ޔ5�8J���Dg����P����r����GK�v����ѣGq�FF�ܶE���.����g�k~���FZ�p"3T;CΩ����ҷ���K��=H���*�9K�N��o���;�"� ��`�5��^�˜*F����'��T/*T��'[�;�S�(��w(6���I^�ݷ.���QvWj�ţP(��'��aul/o�P<��}��Xk�8k�c���&mg!��\�N>� Ng���Q�'�?�ܧ`+�>oߓԝ�2����qu���W�<:�	S��e
������U`(�Xn���י��}񓊝[��zJ�F��`@���28��%�pz8�����ڇ�ᅴ?��-�/�S1�J�&Q�p�a��ȿ�c��pw��̓��
�M�Q�����+�	Pፍ3���1dR*׎�P�iBq��*��C�b�@/�s�R>\���f�9�Ů�Z�	>�����f_��ڃ�x�7�]��x��6KI��V����M��gk��5/��6}���1�Z�Ap�i
:�)�.(��%�WDS�"��9lc�+�bpw�o���i)W9X�-U��$`{����?�:����D#�ve�m���Q]\]��h�3�DP�:��X�}&^()�����y��K��i�W���m�$�7�R�U�5ws�PR`Na�����>�Բ�\���+%����fDN���O��`@�SH���p~NDQq�����q�A_9�F0�������ղ�����h��mع;V%� ��Uyc��37��6:~%!��8YD�#�&�`XI��痏�>!V<���}J�	$� *�/??��AD-�����@j6���lG�/������+G"�K�c�}�0o#�#���ʈ�ZC]+ڌL,�5-`Rkg�n��dS�W��+��8�B`�����#�sy��u�Ԡ2qG��ץ��5�K�Qv��e��Fփ�T�~o4��~/O� 2��:�������a��ݨ��7SDӑ	�ub,��Ƞ���/�\��5i�����p��4$����EZ23�s���W#��8'0�}����W8uu�_򝳣�/��z�����B� ZB	�7���jf��P�H8b�]��5��$��%@2p�G���w�h��=����0O�4a��%}égmm��vh	X�غD&��ZYQ1�����lB�4F���!�T���d!h8�����>��� �����/Brl�͌q��l��z�_{�2� ���29�<T7Z�.�rc1$f���pn�Y�ݢ�3��I�aNo�Vk�x�a�J���
�S�8Ս��f�3 ������Y`1��|}���+`X$��r��ˍ�U��=�`0M}������-s��Rm!��cW��w.�i���o�a��'f7�
�Ke4*E
���Ul;��ѳ~YI����c	�l���ɖ�2�6��)�JN�=��b��J���y@���z*<E ֱ=�>��T���=7����`��r�����^rie�f�o�#�Z��3u����'�F�UE_�׊̸cE�׉��S-� ��qe�ϛ�����t�D� ������_��]��&ֆ6�D^�_\>҆�4/K��t,o�Úϣ���'�o}��l��Y"�����T7FS�ӴT�2G�.)oE.��LȞA�G6/y�:6��� E��o��e�dH�I^@b�ݩ����(/	�2����)I��}�ʧ��ͣ1��I\�F���x�����FG�~�|���3J�P�C����U�d��6J�Tg��OE���V%
�Ʉf���^�|8�~���բ�Jc����/��$�?W��1�&�6d�DRq���zʪT�nЧ�^i����1+�3��@q(T�]N��՗&�����'�A�y�X�1"c��-p�����Fqr���&���1��Ʉ#l��-<���2@�+z]�o���$�fz��;ː���$nT�ވ�'!!�;9���J](O@��k�r�wrl��E`:>�l�vp�S��+6�g��$T._.W��T���[S`�����H��e��`��+����5�~��+.^��P���pA��&���x���e�O0����鮲��R�������dccN:�hWlQ�[hR����� U���Z�n�?~�����ҳ83���[��ڪ���s������h��E�����O���\�7v&Z0B������+�W%@��n㍀sK���ks��) ^6i��
ډb&f��2[����*��f�Џ������ɯ^�֞Z��r������n��FUC�Z���7��l� �w�-�ܡ����& '�3�B��J��2�`�ص��z��J��-���򉟊�j�ˊN��\�Z��7c���S��H�H` է^���T]u"���!�Q�#���L���ʻ�Ds+LG��kd�� �B��
qЅB3H("�k�J`�ac��?^�71kK5��7'��]�MM9��
% ��6;N	�n?{�?��HU�#�J�|��1��2�s��(��Ɔ��'Z9?���^�p�t������.��ѣv�D.lg���jV��7אUu�i1�C�pV����y~kk��Jѡ���}���?Fo빙t��~��?�K XpY�����,ކ��I��˛LI@����A%p�b6N����Z3�!f�"`^8_7\� R�VǪ
���,1}K|��=t���ë��d��9�4g{H�9�_�97��Ƌ��H�W�ۥ�W�i��F��~=�o�m�^����
�rCKOaW��hb|������D�?D*�̿�j�*}��a�����M��3.���}'\-8��kqj���QOO�#NK��1T�e{�c���c�QQ���Y�Q
o�l���C���{ԛ�Ԯh�5\�����H�}����l&aee��4�(-��rm��#�o�rs�dc�NV�)�R[�y��%[�{?�R��3C�ht2�Mi���lI[���fs�p8��u�XO�=\VDä���[9�$�t����LX���̪���3���V\��5M��:����v�����d��o����;�������>��
��cRy!��n�� ĈPC ??̺̮�%
f���>xQ��Ϩ�->Kj�~�nI���M�m���EB�Q(c�#{����	%���U�m/Ӗ�3qd�@7k�d����T��FC_F8/��ٙ���o����\�c<���YQo����8�:��&@%T��m�6@l�1`�>	��E	\��*�bY	ocE��3�Sw����[���u���<�
�m�:n	0�f����"V �%zg�<��Dĩ���No�%�l�K�����/�ݟ��ߍXp�@�G�L~�x�gc�CP�u�ԙ�__~$_���&)}�����n����P�&.f�W+~&��߻v�b�<cP���-[0��t	e̍ ����cmi链��L��B����[ϟ�mu�쯤�(�mB.��ԅyx���(��ܽ{�î|�ծL�-/y�Y��&��ڲ��7���h0b� 3���� ?�lA.���23t�G�ʶ���,��B�Z�����y����&�4X��w�|3��u.z���h���0���.=Ta�J�Ŀm��i��BTg�4���qr�U���QmK�/�+,��>���Rˋ�P��Ɍ�G�L���"��ּ��^i����t4�7%��8��⢋�s�Ғg�oz����E�����T1�'������� ��c��G��22���@M�6�W��&����M�@�bO ;�O�qjM�4��3V���ɘ	���2���MJB:3Uџ�
r��L/^�h�;��������;m�#H�t�װ���HS(Z�<P�{�LH�_���hv�����0Ow�7�P�������Yì�D����D���ۇ����˹���*��	�`UqbA���G��%a4׺�Nef��f��6�K�zG\���ZM=Iou^�K�Q�.�6�u�TRd&�'k����Bت���˟�q�o��X���oe�k�N�x�Tay�E^j5�2�~q4��� ~ߣ��_�s�ʧ�is��D{)�a����:<Bq��������⎬W��W��o�Ɵ8 {祺��d��?�a��/d�z�-z�����%g��_��U��J�̟�(��m��wZD���7ii-�gm�g��)
gq�ӕ��_jc��� �>��M<���tb;���k��n=��LYf}��iy�ɺV�X�g�/�����j�73��ET)�>�d�L��O��gh>)�|^�<�FQ���l
����c��7X!�_F�ĕ�M�E��3�Wmu�Зn�i���,���X�Z$0��{�b�Tm���Z�m;h:�ژ҉F�g�������A���J�T۪���nc��F�(�׊�E*C�-��뛁���	ԞeX������I��>�k_��Q�dAPmˋ�(�_����D6ûc �[8O����T�-1�Av.с)j�������D����Xu+!r�����/�!����j�WZ��Y�͌}s���|y�&e�D�܁��������q�w�g��"��d�3ћY��7By&���j�.��^���.�ϲ%��۪Hp�AA��ٲ�0�|�z�:bM����,c}�������76����E�|����-á��W�����!����5s��vk������:͒d0���\�Q���Ia�8"*�iMs�a�����*���������	m�~�	�
������L���*zH7?O��Z%X?4�ߗ��6�vwEj�쓫����T��V	��2z���|�+G�;` Z����DT����5_�
R�ս�����7�O��˖�Ĝ�8::6&و�{�7·�ۺ�,Z��|r���B�����wD�7n)&��^��Op��)�!=�%��,���m�%׀��=�}�A�s������ ��9l�����/:۠��r��D���O�z��W]r���I�~lmm�)7�*����d(ô��ֲY��7��UQ):��3q�D�kߓ�6i�� 7����>��V�m����r?&���J�D�T��ACf��':�O�i�_�S�tr�dU��T�nb۳;�yXEpn�]$ÏZ��2�t�ǎ$h�C�T�fNy&��I`������Ν{+�����{�5:�:3�N+,��i>sF��	����Ww��U'���'qV���P(Tow7?�~,\�F@εg��+����t�����=; f�Q�c�$j�-7s��چj��?:�nu��3��Iv��i�F�;�������owD}C=�z�{��� =><;�:\Q[����>8|��I���#fg���K���\�@.�|]i���Z���q���b]� Q65��/Fȣ��%���k��R�'^������mi���[8e��J\��\k�y��gO�W�&�P����?��]��m���cwA�6n7����_��=�3��#!�R}�����tD�R�R�H$]�~|�t�p���UV�����z����5z^G?���T�_>Σd��=��=77�}��Z�[}nn�郙tk��R0X�3D�� ^�˛��>])��1ډ��O�Y��(��(3V�n;~�ވ81��(ou�k�2�۸`��my��ㇽ��>^����������������nH�ϙ3S��nRR,��'�Ǝ��E ��YU�����,�U�U=��t�ۻ���s��q7�TҎ�]��/Q ���w�{�^�[jad�9��I �J?�i<N|�m:�^C�cͧ��=��o�`�%倅����������f?�w����<Bn�R���7D�-��0������}�����&
YN�����O��������]��R֯�:A�o��l��J�4��t�����xH>��0�3a������� ��e�����w�%�穀�t����!�;�X�y�1-�y���8f?4��c���/�q��/��E��1�i�����u;Z���K�d��O�9����Y+��;J���a�$���N��0�Y�OZ���u�#��i����ࢺG��?,����bܫʥ�/�a�`��6���XZ#zB��0g<�>}`S3Xf�4V",PL��/��x&��	��&���g�%''��V/")�<R�ߨ��%�\X#�VT���F��;�iV6�_�??,5�2?�9��4{�A�m_�������#�$4���=��/>��!���Z�v�}R4D��3]}�g�V��KB��Ae|��ស����\O�����`>�E/�Y�x߽�{e�� `w�׽��x*hƟþd���y=[���
�=FQ�����:�v�7;��o
�u��i3ؤ���n}�rPVf_4� i����N���2Bc�xccc�|�������4F:Ȭ��(���C#,��3t�Dv����ᎎ��7�I�8�ϳ=�������А.Pc���8������U����O�O]��zߵ"���1t#�5��yR� v�=�����25��l/oV����6�����7�j�޷�鉯ŗI"�2�޼a�~�6I�t#C]�%j��I��Ϲ;P(��m��ˍ�"|.R�@d�+$>����tk�0��=qvC`�<�N(�y����`|}�P�zJ�z.�sS�q!J���I_H|"�H$�C����p��{���]�|6�g$��̳��j�PJ,Vd~ŝ��}��|�:Û(l$W������!V��ԫ���>SbU��#dgl�c�R��q)?�=gI�^me&�j���<V*w͒vhjll4���$�s=�Y�=T2�t�N"��L|	��V�U��@Q���3S�����qX���oQ	#��ʀ�������X�s�	:�m�W�����������þ�Y��:qO�S�_f��i�B���e����d"��(���������$�`*�C
��|�<̓��]�ĵA�7�$e�t�!b����L�tn��)!�#��G]G�yז�c�eZ��*�mO�EV�  �x�����G��.rZ)e�������#�%�v>^�n�
���#�$��˪����"�W�^����v����$�i[OO}���dR�D�;�/l���o[�G8��G	�v��+����h3�t�;3�z�y�\�G�`Q�-}��3̬\I�����n�%ot���@��Qf��W|NRS��������5��\�"q�C���t���
٪nk�����3CY,���w��&�HA�ޗhD{6�B�����կ�p1N3E�j���'%�[J�ğ�Q"��@IXR�wRխ9}��tfNd0h,Z.p�������_��u��ok�H�x���S[��m \%�G�)���qm�|��oy�����lα7�����Nw��e�A���Blu��Z�:�(Y�)�����i;)I�o���xZ(�l	�{|+��w����g�oZ�[�Y۹;��	cٙ��[����`V9N�0@ApGߕ�[��*�|J�v.�#�S�B)�������o$۫>�ڬ(6+}�6ْ��AS��n@PP���[����FG������"�i��K��P���K*;��)E��-v��8K��˛�222D���c��t雔X�7�D�+*z�kz��3(eR�W<���)VA�x_��Ր�g|�/O	�������N�c��(i�-,��#3���#eE>�N�̒��(W���C����5���R���`^R��E�{��m���yep:wB�=2���D��,�� �|�<0����ǫ�z�!�)�k�#���[>���###��G�X�Oɟ<Bga-���<�H7B�*����:�PoC�[�U����������qSTJ.�Z}g�����b�����)1^+..�އ�
��پ!bV��o�P�� k]Jh���]�l����K�S'����E�������$�T�������>(w��z�[��긣�O�}O�S��:��Sf� �#���?��x�8���п�Q��)�.�-��ed�e%%�g/��]b��0�A8��p|5K��זd��F b��+����M�����|�8�<y�ж}��.�ƥ�3��J� ҹ�W���C "��]�\��P������.�渾�1������d�9���5'�qY��~8ݦ��խn�8�V���c5:Q}(r߆�'i��m����x.����x} ]UE�# Ǥ �3u�Q5y��vW��\���cO��
�]u�:��eE�r�w
�5�y/�
�*�C9k�9Z-iP.�C�?��ɢ��[%PlQ�>�4��w����)Kio�y���b��	��z��4���{)e �um-�a�[J+Y4�>���Թ�`3�F=��ݕ����Ύv�焯&�ތ?A��w�����|��ӧJ�m�73��(��R�(�6868ط;
�z}=�%(辪�����~�O��s�ԆU����=��f3~�?��08�Uې���1�Fwh�B�!A����gG^IS�mw��K�B��K_???UUii/	J��J�0�ֶ=�����p[AZ:{�P��n-f�x�(S��(s��������y.�*�Q3�A��9D;�ۘg���*��G��Ⅲ��B������#�~����|�Fe,fh6V��r���,MԝxD���J=���[͡H7> 	z������.6����ʪ'�h4{�����WP���V�r]��"O@�f׹���م�/\����C����'}ܧ=��޽�'�wD�~ٿ��'O���B����%��������V��ƪ�h座k���&@��a:zw�B�#C�_���>#f�M=���3��K�mxG][�]|u���d��ﻰ��KÝ��t��~�?��(����a~D\�c��C菵��݆|u�� C厸�=�9Q�m��x�R�쩖�Q?8
/��<�ꚜ�A��ܗO�p��J|>�)�TA�N����cd0Z����ҫ�}�]����P# ��q�!$��]�����=�����$��>2��p��qY�1��
�y�D�"7hi�+)++��`�jj�>r��R[���0�4}�a�ZB	�D��%��s�P9Ԃ��27��c�
*�O3d�:��E��f���1a?���p\a�]�"9?|JXW��1���}6k�S��n�5���y�=O=Ρ���>�5s&��@'Ѱ�U��������U�̱��Do�/bRo��nͻX�E 5~��a��մ9�eg���K�y�.���Ҵ�S�������(��G|(��UM�[�\dj/A���5�����Y(|�rF���3���:�ܶ<w��GȦ���4ۨRI�βd��^`�����jɧ�~" ��g��2+��me�^5��`x���@d�?ZO+BW�ӒI{Wx�|_WRo���n��VVգAoCqv��A	:puzFD���8pF�5�DIc'�Q�@� ������<c�f���?,cl|�:l�{ܛ1�ǃ���7��@�\3=$+�k�c:��������fz�V��3*��P��i���E|��"�|1�����Jպ�36�e��:����h�O����5���Ik��l!��H*�����
� �����;�����t���j�v͢F�Fcծ�W�^]h)*H�h5���VQ[c�6����1~�<����>���?	99�����>�����_Ⓕ��#��Nː�#Ϳ�n<ZO��[���\�F�I�r^Ͼp�?�����wB�{��)Ӹ��2���k_����q� #Q�>�n>
}�����y��x�u���-(,i��r;1��d�c%��糟���x6�sXZ���R%��p�k��1��'�%��]֨��~<��?16&KT}�5Jm�9 ��jv�6x<C���[���|�r�^�秇v�D\ꄹv�y?��Écn��Z|��W��� �d<�*e������	�qwc@y�+$hf���V����T��5����6I�����D���Y=���j��b����ɴ'�{��Dc��p~���0���ݗ5}�x�b�G�ȶL}t{�k;�A�^�Y��m��L��	Hd�㲒�uMG�-D���M�U���^��]aٓ�˰�=����M��vOd�BjxVJJ�Z���='j�S9��V�����T�.�*�����r�y0G��6���
]Dt��qb�K`?����ۇ�~Ҵe��dCu�Olv&%�>����S��rw>��QR~q{�aj�]�p53C	���^��-3.��}�gS��6V������/�<�]@������zr�x=u
		yu�A�>�5���g�q��4sL���ly'P{�$����b>^�`X~��������4�T����zf�`��/LBL�mv"�R@8V�%��$�4�P����[P�=��8�,��G����������1z:�?XF�l۳^��fw!��=��;[��s���Z��{��'Ƣ-V0����~�j�R�W����S�w�I���ͭ��_�e2�e���2�Wk�#U͖���l!U[U'��� ��Y�\%�1_��_K�8�~��K>�	[9��*�׶��G!�Ln!�a����\�f��n��� R;GF��-�ur�76q��k�?�~Yӟ'������?ɝ,-����g�\[�1��c���m_�ji�!{/�����y���*9�Y��sL�� "3�J��Q��d�l�Twkk+�[ގ�ɝ�bc#�"�\o�?���F�|("��(y����S�_���O�l�mG��͕.YT派3�W�-������d".ߧ����Ȍ�a�;L�j���b�_�64ʡ;.�6�Q��u]�M�"� ��ք'^�g���w���y6�%�+�ZG	���'�,�D��{�k�EC�S恗�ۇ_�s��Dw�QGmjj� ����͡v�"�����O76B��ç�öVFӦ�z�o�B��B��qg��^մk����߲(S.͜d���\a�n��Y���|�䨎:
0�s6^%�A���}�~R}lW����D���m!7x����u�;::��fZ���]��(��𥥥���;�5y�}O�u������M�>���y������60�TR�+������r�Z�z�a����Ԡ	B���}�����}껤����/CP�"�]G�����\����>-�� �/�=Z��:r�D�S��i�%�[��Ɲ�1Ͷ�v�A���2}���ⲲA���np{α�@��B��*��^���<4�w�c㌬��\-%s��#��>� ���yl�� ų�#���Z�
mY/��x����)�.2�����L���ߪ�6^^�S�(��"O�/�~�vkڔ^�ྵZ�eq�K�<� (}��č�Ŭ�Ã�zN%�2Q�����:���?���gf�«� (	;���{oee�W�LM���?��M�M��::�X
���5r��������J���»�f�$�q�c��������'��5o{lnn�������d+�=� ���l�j��A�x֪~�O��`]Gҋ���q�:?�UZ��zи6�~��Z�p���8������/e
�[�zѻ�ͻ�0��i&_b�L$>'��i�L����+�N���ԍH��I&�qo�^Xq��?�oQ�����r'Г�െ�Ý��G����[v7̖�=u�6�j�F<rq��
_�9�?�u�`�����bI���Y�����=�?��D�~��up2��X���vK� ����itD\)~&Ā�����2i�z�
1u.���㉔飰dA�)���Ag�~gv�Q�E�7�S�h�j��V@��XD�޾��	*˫�����>��r:���Χk�E���8zr>m�9~p������n�Q�b��H��"�o#DԢe�?��^��MW\1~�i���X�V�6�b��O'�	�Ķa�n�a����	jrf�R�����x�ݽ	��>s�R�~y�O�I����Y0K�;�\w�viE��'���l,]��ֿ�?w�Bں���: ��%WbLW���D��V�ӌ�\���u�GJ`b�����%6�7~���=�dX�>��'ۑ���d0���-�R6���*�m�M�5�)s�&數nm*d�"� ��gL�4d�{	GQ%�߁����F݌�>T��d�I�jg9C{p=�:�.���)++�5d| 3��x��j�y�Ss�K����2�(:_��͊Bƙ��@\����1������,ti �~2�o��}�\���e��� �<�vD�؀�69��� ��gQeO:���G:�,�=�T��p1D��z���ݾ�џ7US���cǚ��Wc��}-Gm�`������Ɨ����5)��~����47ehO�>�T��v؀8�Cx���0V��'�&|����^��l}7_�z�4�s8�v"�Am�i֕W���}�R�U%�o�!�/�xɰ�K����_��6��ʈ4ڢs2��W[��k��a�2��_j��I�����������Fn�����O>3E�o�s�-�|p�5����=e��S&��,���7���NǱlQR��;	�f	mZ4,����L�.J��;
y��<�N�)����\7���}Ӕa��n��?�?=�ǘ}�M/��x�L%?�bl\����<��3|���L�,��H4��Qr]Z�#���G��/u�4�a�Kq��S8\9?{�O �e?\F.����w 2wdĨcV��`9vU���q?;???~����l�	��q��}�e��o)-�@_��&I(�^cE�@�B�*���3��l���N�v[����`��d��l������i���vbl��P�M�INNND��H��YWǭ���1����I	���gR௑:��� ���E�r�QVFi��LaS##[�ATS��ڒO�;W��ת�4y��=vu-���_�kk�C�H���|�܅z��׸�?q�f������B���Z��H5gu��'�¢�ik=���m��]�%K?�l+��������3^�;��� ��z3Ja������H_�~������+Ȉ���K����
r���7�_���[���qs!�p��)��QQ�._��[�4�IQ��F߾=�fKmB�������O0�;K�w9)�K��w���A�s>�0�!W\ڸ+�V���9/���iX�UZfx�x6���IS5�W����Wx���枙1wI��Ƕ >ܛ �a��N3Y~M�	>,R!x$CΟ�j'�;����h�_���x�G�z��n1�懶7qq��^�d��n����Omخ��5f�.{�p��m���h�L��¨Y�p0�TAY�/zt[|�N�+���N���5nn����d�/u3�����lB��
�(��O�$�5��- b9��3�<�4e��8��SV�|�STøC	�#+�Hr	��I���VGՏ]_ʾ��"�ƫ�s�E�) �6 �����s���ӏ{u>�~�"P�~Y��+@�j��c��ܪ*��<�#9c�Ï�Vʻ��gZN"�;�4���Aِ�R���?���.Ә)���[�7,��H���>J��n�X.��|D#}�"�ӴQ�mKߏ�rz��J�DF=��x���qUXҴ7<\h��:K�Q;��ycor�m\���J��Ӫ� �Ǿ��;�q�=u}}}Y��ubH��m�[Um���y�9`�(�������ڧ2<m�����In�µH�0;�o��(�i���9�E�-Ӄ�J�RAw���I���1�xo�wW�.�M�V8��Ug�E�v|��4R�>�\�/D�'��k���za[zwx�de?`�x�Agc1{�`BrRԢbS�e���5Z�����M���nGA՗]���_�rr0k�������[��*�sPڮ1�?ađ	�å3�|��Xj/ugB3�Ɍ �j�����h�SlL��u�D���ҿdk���q��Z����������9�Btr#n�ro�$��{P�F6"�3������4w�Gq����vb*I������먁�F]�I�ۍ;��k�l���'}��ތ�>�~h����dS��IѠ,�2
�O�'m\9Zّ*NP�� b�ו�`���~��# ?4�C[�qe�^'DƠi�p�h�\�� �-g�>_A���W�/���b����>���.�NݍtP�=����f�T�Ue#|��*;g��`�q����c��e�]U��]�l�,|V6b��QWJ��!��MY����Y:�ʅ�8�}BZT���+ߧ�$L;���Q��g��O��x��D���1ɗ�4YdF�Ȯ&Ovk����@���QJ!���'�Q)
g�ɗ�-Ǯ<y�v����O�d�����ã�LGz��_R*t�wZβ�r�s���D3�x�&���s�0���<Ww���&�}���ri��'G���ǳ5e��h<���Hh��t�6��{X���>�/6�.G^�x���L2�cs��2x5�`p�E�e�	��`�1j<Z����.��?b��j�^��,��|�̱���~�!��f�P!���?|a%��[CzZ�g�!7��-q��p���Cȫ��Z\�)�����2n�b��Ms	s��,C�!��A�Dn���@�R}�kY�@�g��@Ӽ|��	 �9����Af��g�g���2^3ٮp-���"�2���������M��kU�o-���ZQ��G�x�2�_�zeXx"E@����b]���g�/ީ�6iQO�6	1��a���G(����$��=Z����0����+)!Q�D��S�K�r0Wq3�����~2������һ(r�~���i�#���F-���� �'���io��e#;�K�^���q�~����aoOw�@��"�-��-~ߟ�i�.�>�\����.A��YbՓ��h9�ꢾ}�?LjI�y係U❝X�"2XdI,M��++'�J���Q�)ZܱOh���s����2@c��J;_GG��~�/�?5�Ca�+(�
 �������Yt��I|�"�R�s��Ѯ�x��� �ʈ�3��e줒�H��������.� Эtu�hϏۗ?���C#W'�H�;6g��Ls��>�^�kF�O<7{��>7y,�2%E&�L��I���Pa^�&���hoFC��*�J������b_��i�j����=9���}���}�����\X���Q;%k1נ��?����+hlT 0�����8�R�LY_p{ʇn�@
?�w���ߛ�l���?��z�<�����d�*� 4�K�Y ����nH�Rkt=)����L�2�>���@����q�m���SZbwY�i���e8����s����h�R�	�
4B�p�����y���,߳��;��o�:�_~���?���ÀZ��m<M#q�8r ����#4� ��w���4�vLФ
&���=S�-�ܻBC B�ջ�����d`bL}t�l��՚��Q��9%�S��Ĩw���k`.�ML43'��f��v�ku��b�Ұ9bFm�pm�6���@�n�+Mp�E�A����&���m�JG>���3����(���_�s�xx?qJ�6��@�ι����'�!W��D�1�e��{E�1߲�J�7���X��4/�_oD��!�Tr8���v�>����ADF}Xǥ����h߼�e|IIJJ�S�,v`@����pK��L���c�b���'x���H�S�I�把���a��Ƿз�M��1:�VQQa�E]���4}���U]���36r�ܺy�i��3Zr�_}�>d�,m�o*\،
�������^��������Z�v�!��:`݆^��vȻ�AA�j�����(F���ƺ[��f���J�3f�2��������/3q�����{���������i���D@��	U谡��Q�Z��5Q�u^�f�
�5At{]�AP�z���1����;nh`�S?)�ޛ��͹��K��4�v���N�y��c�����7����?m�44o޼�&���V�����}�Ef������d^�]��Yd<�;�f��y`�Wĵ]�[۩���_�B�b�tS�2+-my�\��&""by�;M>O��q�;~5���Y�;JJͦ�ƲQ7���ׯ�H]P���Jn�\Z��������w�-���B�ދ\+tE̗/���@�1��A��nRf��m��7
��ꥂ4�}��l��+j 0�snr�_�����6�<�����ihe�ˣ�h��ԏe�9�]���6H�uЇB��@��h�ף9��z�}�D�F{V�2���1�w;S�j
/)��5�¾a'h�F\�k�3�W��.���$�d���8��ņ0s�_
�x����E���������r��A�K0����]��Sl~���5ж^'�l$B��2���������A���;��X�v}��X��Q�؜���5/9�rQ��E��;���ʾDЫ��k��,]��u�y��h�!KW�&��at�{H"z��S�s4��N���ghN=tr�܍R�N�N(>_�?H���~��X�����Ms���Nq�bP0a��q�љ.�����ODd ��k��]}�q^Sݧ�pHU�+�|e��az��:? �w�|��ҙ�*�ss�*��)c�@h�v�te�:���>V��3B��ji�i0=�RsI����y]��UK.�U/���y������������-y3&glK-�3"�D��{�� m6�X�����Ų�������p"v�،X=�A>�[��R�L�<����j+�;V�K^4{�x������U�_�l�at�^U6�7��$�M"n�����O��J�oq8�*��_��,O�jwq�/��@�ܒȧV��ukm��mJ:\o^�j�Ϡ��z�:/��0���=ݷ�S������iZ΋���TO"n](��&>�]Z�rK�`��>�E���r���斲�h���i�����<�[F����OQZ[屎�$�,��Qͷ��"���h�|�����H�F�k�,��'��E��9杶�tP�5gD%�ؗ�R�7�{cs��~�氃�b3�͕Q��v� �5���ǡ�6�%�(�����uE�C��P�[��=ȫ;��C��.>�5s^�� j�����\Z+����|�3��|����ӨtJ��A�0�)(�jZ�8�e�O�-���3�V��kp�̵�&Z_�,�!jl��q hg6J2�p�����u{!�n���%C�Œ?���ۏ IIF�lo�,X��I��$#��9�07ƙ����궞�P�>^{p�j��(�摷wٴ����p�W���ϘS�I_�T��)�:cQ�2�tt���B�tGZZ�����D��G��t-%��7$���,�A��5�a��i���AAv����e�C�1N�*�
���2���o_�,h\�����=;·m�#�%)�.5�h�r���96#���XAkJ�n��ᚔ��S_����cٝ����x���4�]��6��%w�`y��l�Zi�a�/s�_���h�Y���{��ko�z���\�v�!���Ehy��C����3X�����v�P��B\֢�;ލvX-��ğٴ����������X!�O!xki�j�B���x�=ۤ����t�����Nc��u�:bRV��}~���:i�*����m�U)�I��ﻷ�-���K{���1���і�*uk6�0C{gi���5F����k7�����!F�$�|h�wY��A��X��������o]	n\_>��}�Z��7ۻ�� ���x"
��������y�}��o�8�dME�\G��BOj�=�H@�O�pG_�E�ܼ�2Y��=�*����޾�p��jUD=��D��ͨf2.5eZ�ר�g�EK�w���xg�j7�aw�Ҟ5J5�,F�_�i;�+6+?	��'*B�]�t��Y�G��%^�(VA��;g��3�H�v���
�����������ؚ��/~8-n�0#�V���"�y��
B�1��ġ8џ�	I���'qۂh.N�kW��°�U1DS��G�C=���_NT�@�:/O�.<Xn߽��%c�p@}&�-�)��5�ih�����i��[�aV�{bo��\�$v]X8��\Þ*��O=~٢=W�Ɏ�����5i\S���I3��4��&�v��jG��!�y��{�X����i�ۤ����L�Pch[�=��2����WE�p��:��h���xU�a�3�6�[v�]z\q�l�F�v�W��2�joN>P�(�@��u���F1�߱���K�a�_��G�~�؀��7�%��S�2^k ��q)���\�#�p?���,�+�mKA����5Y�����2+C�$~�����
zx�;�����@�$��?�&E:�W�<[I���"I�C�8���_��g��%@n
�e�����%��{�x��C[:���.��(�dJ��&Q�+��9A�ˆ�a_�\t4l9�!Zr.z$(����r��1��(���gH_W�y>ڥ�p��Y���WYT�T��Q�1�T�V^s�%(i�Ä��l;a"�B���G�����k�zF̈́��OgH��7���
<�����:I�G<��$|"�ۉ��W����՝XyM]]jfrz(���.�Ko��UI�?���\�A��U��N�ok���]�$�ݏa�gm:E������_6��Ƃ��4��E���:]��� <��\6>�;�>$ %��34���&���˂���}O�C_�d�͢�^��ٰ+	����Ҟ�n��_�b�V4�����=�ʴ۹�:2#�Y�$
Y~+��0]�!�׳V�KMM� ݼ�=:�ִЗI�zdI��Q�a�X�k��?�3�_1��.�]�V��>�x5Ӵ碦�<D����EEK���KT#�$��Tq�ӧOÇM9��+���_�x���4=-��t����q�uú[��q��u�7;�������_]��:���A�-#�v\V���鸌Of���.������D��sɻ_��z�pV�34ߙ(lV�9�@*��e�$�g��H��T!�wxxP_� [�jJ�yW�����L��8
[6Ԭ�e&���H����|�� /o��~��Q��g��5i���,LS(���PLLLUЦ��<�Ơ�����VjŚ�����rb���^2����Ю�>��8�`@`���m���K���5:��\����J����-��pC�V�L&o�_�:�;;�kMS1a�i@5iJ����l7�I ��9df���ozΓ
�t�#��q��3�������*	1e����@ar,�5[^]|�5l_x��	���;��q�V��q"�f1�/����AYȫ$c9�n5΄L�a]�P�˼�2�UN�Y����,���cGwq�1�L�@��2�so�R3x�O�Ձ�x�����u�ly�07�`�@Yk�Xj�,�[ʭ� �4;�][������b���=V�M��
X��]M��c1u��A<�ù���Ym����+�?e��/�."�W=�o�4'�ko��$.��
Fěs#�kB��L#�2�\&�v��e�W=���s��ЉeY��_JzN�S����u��+���h������<Vq�g���F'e��{�j���+�����DY��˄)�L+�5�b�jw���T��o�n��m�6j�!�v�G.�_��;�|�u]��M?1s�Gmw�1�Q��ZUdN\.�f�E�Q��-sR��n>*�ޘ8;;�b������}�ΰ�i��2`�46�[�p���]�j�U�86MeG\�C�����ll���)OLL�ұ�{��۷i��F��	��k[.�**/=�v� �9�����7\/,���R�R!hC�Ĳq�Y��p���gú��6�M�� �8��,Ǵ� t����(�{���p��ݢ�C?�l�?i0�r)��;��!�N75*��F�~p�2R�
�ן;��>﫣}�)Yj�q���t�Ů%帷��t��va>�)&���:~�yK���wn_�ý������1	���j�;QdN�؄<k �^�a@�]r:�T�k�Y�#�vdn�<i#�8=b�o����n��g�K}2I��pKc���e����[&��{D1m}�z�a�� �"��rW{�$��IC@�&��/_��K�ޕp蹪��7����n�>|����L2z���m�5`�k̳L^)U��?��Г�qe�m2�ܛ&X�]CU�;�s���($���6BN�X�i�X��>o/'vp�O���&#��qvv6_?
V{��	`���ܒxn%˒��:���w�K�$)l����En���*��G��7��?�_#�e��P5��U(��Z��mRq�G�;t�qD��|�m���_�mG]�YX�m�p� �b��OxZ�����=��0)w2'\C/�����c�Q�rYgư"õйV����8f�f���W��a�:����J)��A��Rc��.�e_
K��߇�p%T������-����X�M�b�4��e��"��4{���	�|�)ڼ؏T0�
�L�`6��_�}�����}=�딄,����rr_�Qe[�^p�Ģ��jg׃3���@E��NSKH���6�����z%]��ʷ����{�Ii�EHZ[?+�����r W3ʷbD�4�M+��5�f)���pIp�C����V& j�˃`7Xj�J��}��-�Ƥ�4��ٳ��qOb�ܚBĢ��
3s��}0v��l�WG'�̅�3� փC��O���G+r���6C��:;;��~�~�H$H��q�{��>=��5Z}k�j'�NPA~�L�FImvK�@�W���M����~['H�x%�PJ��N�3��QB�����^"����*�+i�&f�m.����~�b�;p�W9A���tDGA�P^I��e�g7ɻ�xG�LTM���_:����p��ͯo{����G�~%�'���~��Y���k��������{���78-W�y�D)��㿧X�esU2�a;F�q-i���q5����_Xz���Ų��ƭ����a***6_�igȔ��+�^}��������o�����N�ھ��a����8���g>���r��Y%u����J��kdj��}Rb⧆�_����9�"D���^L����_�
aMӇ[X�m?�jY��<�� �BFGG������_ ,��x;p�b�ud��eU�)!H��D��>/��
N}T�q�#������ͺ<voBr"�g��HE�7��J�_�n�co'p�No�C��Tº��Ty�G�qk�&�=���!�]a^���CbJ��=Z!
m�62d<ng���;�mz`��ފ��BBC �t�$���?���z���B�(��vK����	ZsP?�҈3��$�{XouI8�Lk��������q0�;:��>� H2VaXh�7�=�>��%�X���X�b<�0�lP=���M�{��;P��-��t���w%n֐��+,���Zj�0璭ru�ȟݩ����i~�\�d?�z��j�c��y���P����λ��'�Τ{	��¢BCl)؛L;s^u�;w�S�uP*�
d!��]f')�^���.]�9X�`��]�j	Z��j��R�BN/Q��4It"�Y��a�������s�5���6�AY�"��JM���(	5�v[w�}󾩦sWnX[mv���w���zEdP�^b�:o5<[^>������m�#Hj0+����j�V�d�{��oB�^L�(��뒁 �m��t���(:���e��?K�{��ZR��;�\df�B�!n�X8}�=ش�l�9�7���F�˫��&V��%	?q�趚��S��F�3����J߾���L�{e�� II-�������L��σw��\�M��S�C�{ �(�xnz�2�<����t�-P��X���Os�־�޷�w�$��o@�)lbh�n{�����,�E���ݔ����9��&��w���'�Cl|>hm9ԡj�<&48^S��n.�	w�U���4�_B�F�;6HBmO�l�6���L�CNd��k����i�;�÷eW����c�SÜ9���,�?\���������� f�`�c��멆��v8.�s���T��Y����y�y�hӎ�j��z�EM��}��#��h��ߨ����B�@���5A�O�G,���,j�Z��'}���iK�J����-�3I��bwC�p�����\�W��KT�6���حV�f$B��{�aq�l��
��1�q<In1r$�JzS/���֎X���p$�@J��<.����r�x��0�U�q�e1 u)
�j1,�a�� �?��B(����㼝��c�
��n�2��ݣ)�#|OV�H@&�|'9	�Z}�گ��!�A!��=*_�����y ~�����
�����U�w%<H���~+)Z�@�1sss�ׇ�>�唫^٫#b2d��򁭭m�H�ء�C^Z:1�����k�gG��"A*��x�D�[#7ܻӖ�Ը¹���/�ѯ%���*)���Ltd��M���o��̉-��i��a�(�S4D��:����rY�ypxH����m��n��� �[ҕK6�����b�A����+�s��3i}�����x� �C���������'m�Q�������VT��e�.�1b�iX��`�Qlu��snWp�<2%%��2��~ �����ʉ552�u�.�_R �<X��Z_��5��l�G�
�Î3�i���ϧ��Q]�>��VVJįRݣA���O>�}A�o��
��c~/)Z�(�RWG*Q�=0������ۑ�j�A��r�C(�[�ѭ6i,����PH�n믔���e��o�)�_�W��@�eNXA!�\;LH�{H��5Mi�DEKc���|�2��[�K������'�q&����YCGF�.n�KVJ�r�M@�e ���^P$���UY�*��n�z���͋�"z��U�&tΔ,�Ƨ^��qN��{ ��P�~�}7�ųN޺���b3i��e>�uB.ۥ˗'G�����`�Q��Q��j�$b�`��9��J�T��w:��U�^��o�~?��A!x�i�=v��ԆtI��yP�*����5� k�v��%�F�a��d*�ލ��(5`��n+5�sC�i��\���p XS����y<^�	�@��}\�[��يNw��+"jW}���^kj4�Ii��n#Ä{^���ݰ%���Lb�G��~��Y�TAK8��X�6.^�n<w��5nYKP
�jZ�Uc�w�f�X$���׌A��w�j���"���]���ه~�Pd���,�_l§�VW	3]��s���CH3}fh�6��3��Q���A	��ٞ����;ۦo�ͪ�Z�.P
��ߩ�m1�����Q�˃��wy�s�6w�0���i�4��B1���`{��=�����YX��]��H���0Tc�vA�>�u:xM�K�1��K�ԛ<�w��Pݫ���[� �r7�]ag/��S���+ Z+A�����
��̾K`���a��ע�����_�h�FԮ��>��Z�5�1�?�ʛ~���Y���*Ȍ ?����G�)ҧW���"�CL&��99~_�W	�hf�����2ܘs��A�����g6�q�^g�a�oG��� ����������\�M��[��k�\{ioܸ�[MZ����^]��~>��ߟ�R�:'tKkj���A��:T�D���a���O�G󁟚F}�ǐs�Ƃ8Df��D�w���}�ק�Y�jQ�����8�sg�bj�0%4�͹��{��S!)kY���^"0��mm^�8x��f?�_� ���M}q���H"�ۦu��YV�w��Y��(P/�V���!�UӢ�Y��D9/y)p�������KU��@��z`p����CW�o� �8�'f����vH�,<B�l����b�e��BS�A��l�/ Z���ɠث`���-PoYf1~5�u��v7�w�QX����e���z�E�T��:�l2k�I���8.��-�����;��, $pX�F���6t10a��c!�����bl�&״��zV���1+�X��M �F8�.�$�4��� :��
�9���6�zy!U��c4M�'Z�4�Z�tڇ���,fh_h��~9�`��б���F�h=�[�=l΂��U����E��*��|� 4�^��f��e~Y%C�ݮ�O�<��F����B�9��ξ>�$)����Twۚӻ7��L�k=	��%��g	�x��P���޶)�H�V=�C��f1t��c�aM�♝���D��d��t��P"KU0r�/��̽>�6�pЮrM�t�����x���8yr�S�Jo@�����o�җ��:qc��sD؉wP���jOJs�uo������Y}��]f>���?s�?���P�l��T�3����L?$1cvΖ��L"���!�ȴ`7��u�����/�{�w��LQ�Pk��w���Z��M6�w�����Ϗ���\�c;��"�t���vO%�͠ 7�R[�9t��q ���L(��ٚ|�ޣ{��^53�R��7��Lc1
�������~��Wq��nT��O�^��r���d?��/a�Ш+�$�5�fJ�`��|�i��FU�}��acu4���d����(��c9C�@��Y��ӯI���paV�9��p��}S?ā
E7�y����ޟw����-�PD���?��6;���Y
2}Q��;�V0_���+����ER��Zp}V<h��҅��.�of�x��cB��cկyQ��Q˥�%3%��ȉ������ia��ɗ'�*kM���9�CNQT���: D�5�	���'xܧxع�e�?����cL���G�O���	�~�u�4�U���J�o~��H�1X�j*kI��\�Z���E��m
�@�w�à�Jꣴ�m�fc�/h��UJ�����m1��}�%+'gV�Zn�ޒtZ�,~�����5a#�w/��j�\;7��S��<g�˛��2��� J�@��.t�O2������Vf�_ �_�+�8F2��<h����ѝ�}���y��/֠&ǘh��;^���k==����-0���X,�x�GG���fC@F�M�@ 
�[ao�|�����^Οd`mm��@�b��1Rlm6����UUv�t�+�1]EqéŢ���%Ko�O5
K��l��{<���eX�svC�ٗ�\!q��3����u��q�	�ٹy�}ו���Qǽ}r�pQޞ�$��Ey�kQ�����u_��)���
��������Bj� �����xc���;y��ז�H�,BO>P��Vd&a�/���_��G��Y��a)4@\�|�Nx����a4�C5/�������4^��Ͱ�`혘}���>R�uD��0��B�������<M�zdT�}$��6x�F~�$_VyM�ud�z�cpo�XXi��ƳgƬ���.PP@���QX���{�^Y��i�2E�X�kh_;�Y�90��;�G�5�AH�O[�j�u_T�g�")Uf���ԇ��QL�����[bڃ��Gb~�����¸��]@H�-�Ǘ�~32�
�$ʔ���T!������;��u55����\S2��#�����ZGD]=R�`C���Ѭ.^��-aӼA�+���D�]���?g{�`v�[]4�����Yp���`�(�EWtV��T8��Z�����r�&L=�N���jd���Bҏ4���͹�99���Z�źUJ-ӓ�P(ek8[-&)!�#�����,��%�ӡ�&&&{� ��1?���OkӒ��x��.C��ˈ�N
C0_�/��������w!���U:�}uU�G����Y/g"���GjVʻ�J��Հ��^��z��T#�!�*�1�X�j�Q:T��U���r 
g�Sm1�[���U�!#�B�c�"��3�~T�Tv���Z��?�����˃�����:jE�_@ ��}�bc-Y���}d�y����K{�U�(���/�/�*�n� �@�׷�T�ƻ���${��!5�dk��@o�B��ز�ti���\#�w��=��-����A 9���V�l��w/l��[[�}jpc�����p����bW�������Ћ�����e{�huC5��;�e~�Ei�w�`��Hm�2�ga��ḭ���o1����\X��"\$��#$4��⭗g�7~�2[^І�+1?)a��I���V&%��,0�פ6��~?�\�F�� �T�0�@ ,X0@\,C7�ɂ���#���< ��F��=�������:�h�����/ɸ큫V�UG��A�&�֢���T�}UX���I��@~�<���zs.*劣���ZY	����gg��6�x���o߾U�%���ddd<E�i��[��H�'�^�B�΃s�ϟ�1�;ZdR�����qr�S�eG�o�n�����H�_~�7�ۻ�2d]�S1��j��rӉ9�� f�1d2�� 	$-��ؤB�?}q�����u�����l�1
\b��|>�ཱྀ��^U�i�A�����;�C�����xȡ��ag����֠�݋��H1V�\��_Mg�Մ�����26���P��Lp���
=�Թ��~���E��3�;tw@}�S��}^YDO�Šso�c�9s����-�r��U{GI���D%f*l[|iL>OO?���ĳyMa�:��0J��$뫊kl�U#}++����P�TŲ����S�X-P�_W������Z�~�զ�9����Ԗ���[�r��3�T�۲{K-@�I]W.4�B-KC�h�B�p���{�[��� ���=��|�9�{N��je	u���2"8�aW�,�a�<��\�9ދ��4�4��X��o�Qy��ɯ**N@�#"jVys�_G��̹�yC�a��/�I}�0"�62��k>��3�/�튟�lth�b?�=�S��L�C�|��I��o�f�6����8팡���)��s7���F��W��-%����7+�	�ޝ�Z��N[�^(G3����(�-~ۈXa'�^�Y��8�c��X���.�oxuU_ߊ)A�c�F����߼s��d��YRT��B������'ܬr6�5�^�u�P�#M�[f�l�����H�H�!��_�*V"������OU�sE0�7���~��1�͌u*2�v^�綸��k%�>8Fv���D���'�͉Swd"Q�_e\���/_��U p �^�������"v��%f
}�13=��X��X9G$f.//�"D;z��g�`-�>�\jl@Wf��?�:� \���n�ѿ��ry��V�P)2�@ !�P��8�|OT�ʙ$�䤑�?�w-ޒ��(��{?�]j��=��V]K+������h�¹�y �a���˱��t[��z�`��TD�)}ɺD6A`ק]�@��z��i�V�0a� ��A������R�"�^M���Q�G���N{v��u��'��졸���Q2s�q{��o�j[P |�z�f,	�Yl̀l�t���ֽmh�mX��/R��K!  :߭�+�Q��#��8y��ػ}�7˜F}��~���TS��V�89 !T?A�����T&�I�FX%$$���аP,���D�fpJo�-]E��7������UhJB?�2����(RmF!!<�gA���Ξ���2�y��Ff�$��	 O�H {M�,��_�Wb��{�1;՝-l(��'����e�x!˖V�i?�W�pvQ]Tvܽ�bc�n#�6񈬬,dg:�fP��dx��j�+�Y��%p���>|yY���T:	�ݣ!�{�҆�*{*�73���<���$���m?C�����Cj�{���(Y�0�U:�+<	ׅ�b��e>U�H���Lr3��f�$h��3�ѓ@@��b�����a%x��+�<��>��YK?�XJ�;� 3Dz���dF#�5Ǹ���D�q#EW9$���\3����}X[�'���*�� QI	9��0�����(Y�^�>_�6��.vA
����N ��)l U��K,|}s ���>�Y]���F�Ǔ��E_VRQ!!O��X�˩�,�uo���r?�s¾�GS�YD����%��T�����#H�����9�f�p���6_gGw^}r5����x>chP�I�A+BV�}r_KKK7=�/!o��B��TGZ�c�>�sJJ��t5�g ���5*�da �$��J*F�Z߾]����6������ᦩ(~G�E�J���۽�w�,��/�5!#<ϡ�d�`�}�}�����_q�HM�d趶;��켁Y]��5WG��a��Vܛ�0���]%X��թ͉�c)-���9��D��0+����hI�]uO��w��<z�@�:�]Y�ƥSc�S9�{��(��w��p,y0���5��=�D���Ml[\%�Viz�@�u�w 쌆ïݒ��nҠ�'v��AHH�����7<�C,Ь��[��Ug�)w~^�L�"��C�XE�)��@`À�;7
_4��B{ȥ��Α�P��	��� +� V@��*��0��#6� �:������'�$[�K�n�=��}t믩�]QGC���F����-�#Ǐ[Y/9"R�����8Xx�^�?s�S��ۭ��ʛ	�5 ������� ͢���MU���U�����̓�7 ��.}z�&ڴNa����N?wʄ�/(i�4i��,�k݄��E��>}�}['c�<,d�f�jK�{-q��V���>�zC̵?��:�����h'j�fy��' [��׽��rj�b��ri�E��"Pghg
��&�KB;�e��@�[3#c�������\���75)��@_benؗطB��|N`�ǵ�$��JT_/�/���"|	�ܤ��<U=W��e�m7��砠 ���t�r�"�frcL�
��>���f�Z���jy��~�Q�Щ��܆�hW�!@�;3��$N~��}v�0���.2���P�zw���;�]��-SS6�n��ʦ.��3�Q[@w��<��יL �հ/<w�� �\�YG�Da'�J���+�K3�ev�r(����t(ޗ�*i��TH0K҆�?�S�����,˂o�sє���},����%��݂����o��}�[9��6lТtL�CA�co�e���r��"�T�"6�� �u
�O�p~��uK��ajx(PS�g�-���7Y3��$���\>bX�:�w�.��C��L��p[[�K8G�`�(t*����ߎ"�ͯ �
�ˏ9��������T��L�E��b�?��XJ��?�l��M;*1�M���}��<��Y�ַ��	!�����L�,�����,M4BS �d�:	-���\������9B���4з\�ZJ�bx1�Ηy:�����~w���>��n���b6iOi�ٽi���q��l�B䖝rW2/u �,�j�Ң�b]������ �6
��̙3��o}%>]�������o�ligr�G�7�Bm6ا^<z�/A�ޡ���/���Xn��-LVv���¹s�M�?� �@�?ck`nu�IWn�����{�yi���'���-�B>7��p�qi�E�˰Q�8D��n�Cٞ_nR�(vO�	B�.l)�GJHV �/�Ȟ��5�J�"X�/�>��Y�@�mo�����F���N�����]H�o]:��N筌�)����*��J$�3�߫��k�cqS}��q
���>��V�f�Uk��"b��/����[�I�gy�+���QY���A�e�xW	�ۦm%ld�:<�(}�e�)N 02��YY���D� 
�ǶV��8��φ/�t<ٯ]��8�;WB���l�9j5hr��r�(�̪8#�dO-jo�����L���6Y�$�*P�~�5��������'�`�> P�&B�@�ono����*��|�%�OWu������W$��{�l�l���*�J�*��K[^^6�yh޾����`V+꧔�d������Q��JT�U�\W��l��Dix�O"l�)e_h����{�� ����d1��t������������Q���$������O+��;�I�����w
2/�?��6�PaP�kI!�]��pyMX˻z�g8�ߥ3BL�	��_^��`��]�(��Fy�4�h#5��娮�4y�k��n�+ݨλ���u�O���Z��;�'2�:���x%�������N']6����~�[
Q�s�h�XpY�A[�Bq���a�B��E���	36�k��<�>�X�
-=��`���Y�E��Ȋye�Nxp��H2�l��FJ1�a&;8<s�����[�&E3��Т�kut�4�y��޶��2��(��(��I}0gz��h�z����|�b�I~�7fʵ�b���9|˷�b�$�{g��iqi�.�Z�5��<�g������/�X��_{�,R��o~{���� ��ԩy�������}��di�6���{���I#X+^U�;K��4a�EX�����y���ËJ��.���&�6E�#"#wh%��]obo���&}�\n^x�cc�����R�f���$S� NɴF̀��E�(U�⍛������4����5h�9eB#�)�Q	Xc�x4z���VS�H�^����3`�E����du����$���z+������z{Ռ��\{��m����V�\f��Mx�:!/ypyˌ��T(���}��)	�C��&�����G|�nLP�ŮMD1%sK>]�;�#��W�����u/6�p�XZ�X�=})#�<2�'f<}��߽�$�:]0&M%���2��/cFti5���T�i����p� �Z++����u��@Z:|s�T��ru3��p��"*��:�z���X���`0�_���$�f%�ʻ���O��'�㆗�:ci&�mo-!p��'�[��7�nm�g��V)'�J�����,�K��e���r
�W�4ϥv ������A���_L����@
�h���JBߌ�����Q��T���k ܿhĊ�T���e�s�D1��w<U�wu�Aڐo~
U���kU�+�i�G�������V��wH�5+��� ��T�v6���8�I�k�K��P	J���� �������ρ�<�8[\�E�ߣ%��C��FYra�,:�	94���b.�MG�[LЗ�O��t��?UmPno�c$
�:��榥c�2���:�1�ָ�:w2��C��Rxı;y��vݎ��W=~l��a�F�L��$�z�NY��qC<q��G'e�H�/���8����Am�9k�`�̏?��-2j�����z���L��CP
E��=�·Z�5��q���sUX�����f8������I�-]���]���;��a,�(=�1������4�Jw���n�ю���:�v�c:���r�Q��#�7�C��,��K�4�4S��~�:��1�ֹ��ڞ��-+����Ą��f�i��oq~���&���Qv8�P�%3f�A�JJ�ޑ&��$���5�KG�@�?��-Z`A-�zG3Q���m)��rɕ)W��R�(�CH8%Xà\���:QN$�-K�H�uC�܀��xp<&hbj�^f��N��RL��#�z���~di?,����x'X���_�!G|��і�q�NL�IaT�\�I{���ۑ2���Q��[��(��}j-�`���o��A�y���w�~?Mb(��X�VzL�$����c��zkj���� j����'���?��6��ŝ��~Z���+8�=xȣ�ļIX��E����g�l�r��9�Y�>�
ɑ	*������^�+��=�
�>�MM�=�	���{�Z�P7i��4<����ଯ� ����m��+��cT3�㏡���������6�Hv���T��]�S��p�K��r ���8���8'C?�sBe��-���8I�j��V��\	������ޝ�)�@��W�p<�"�tb�v��[�Jc�"�a��b�?A�ף��#�_�%x����D�fE]�,�������yd
�3��/�7�e�.�s�6�-ޔ)
�5�8G9�v��PK   �}XP��/�  ǽ  /   images/f42d805d-3c79-4d19-85d7-77e6ec425ca7.png\�T����"  "%�R"��%�]�J7�ҝRҭtww�tI���<��]wݽ�Y.����;o<����U�GA�C���A��Q���u��y���s}X��y�($����������H����,{;)�z0�VP,~gN��,khm�l*S�6f��}D!3ܤ��VR�q{�Y\ÑV�]'A���fӵ4�ϓ��q�K����y���q�=~<I�����ӗ!hG{��%�M?�ă���w-&O���;z+8��Q���f���~O�&��D���?��e�yJ�@�-B�����z%1�����>&]���b��bp��W�	�H(a�o��d��-���Q�+4�R\�xWe���*.4�����oq�`��F8��c�L{p��ڢ��}
sR��z�S�!�����w�
^~&�*]��R�\H��sݐq�g�A�*�{��p���_���tcd�=㬖T[`��e�b�^Y0>Y��҆�R�L���y��up������$:�+􇇇�q2o��h�ۮ|�6 +ݐ����%T��0+�U����"���7��\��A����'��KF�R���������Jy ��a��υ�;�f��J;��	}|��j�b�i�]�|$1�\��s� i��~b�ͤ=,
�Ȁ��I>��[$�m��-"�c�V��g�~���'�����K��k>:,��.�"C����H��3�_$2^.<�U��)�	W����
ٟ?���*ȥI��+̕b����b�
�Tm&��J�](H��7{���w�xc��%"ҽ�Q�Ύ���<���Ͳ��kNtttfף%���qj�ES���.���8��a���A�Oԧ	�XH�?�����K���s� ȸ4w0��.��\�g�?��涉�Ȃ�E�L��/ڿ�q��1�w�0��ßj0�������@*����8�����E{gm�R���AY%ߣ���<,�QO}�o���04��=����_/��W��"BB�N�l��0�\@0~�h�U&H$�=��?�W��� u���YLAL$��Sh�,�٩�ha4b>�<P%oɁ�@����S����ez�R��M�/6��C�i.f�����oӳ�������S�ae*���r�|%�|%�MV��0"u�T����B�l���2w�$����u?I.�ꟆU�nn80�����00x��0�������CnbȚ	3y�6��7P�_,��
D*��{y��?�%���&PRVN�!��d-O��6�_d�����ѫD��,��V��c�݃�k˩�$^����96�
Ll_Q��z���)�����%��'.�7�ٓ����>�$g�_�1vm����
	B�^��z�t	
��;"$��UU����.���f�B�փ.��'�����뙓 �vHOW��3� ��S/
�����?vW7��KF<jF��Z�G��p�����V��GF�;�uu-7K�Ɉ�(!�a]�"���T�OM��<7�DE�待6���V�!�iJ�%9�f��f�����S�?2ޤ��CNS��m��^�?=�b��vjwZe����R>(���/�%�SF�'�g��a��渶�0n�C6�l���_����o���ͽX"%ُ�
����cka��,x�|t�|rE)Q���;��Ի�I��_[���W1Նp���eK�w5���b��k!0TW;O�/:"��M���{c�;�_�|E$��E���+�eE���K�k6��	+7�-��I�t�S
�^�r#^���Hw�k�����!��#�#�k�K%%�<\����D-���M�=	�F�dq�8�455[|�$��42�˖�p���c�٢Q��X^E��\�:��祺���Ĩ�sh��7n���sj���i(2T�E*aY���;�����LoD�Ă��G�����=S'owk���K-x_����>I�����D���Z���Ͽj9��!CO�7���{�K���dvu�o�W��aA�sbaqS)�1K�"�w�Q�ӳ���,}9*�΀���4[(���8��`��}�慀!.�?�XT==��0�*T6Ư�"�ڃΏ[���l%E�R'fH�p���E�� 4a������ײ�|�b1�c����aID��9wf��X��Ku�0���d�0��,^�c?_*��+l"�.�������k���Թ����ܽG
u.6%��M���
br��O$�N�?�?�bi���ܛ�\~�u1t`�0�AS=���~��3��e>z�����������uR�@�h�|Y�+�9�qM47��B���F8��&��O���\�p�}����uJ�y�H�k82z��_��9�"�5��`-��|&r�LS�Q��+%BŠrV,*����#om�.ל� W,�}9�@�p�H�����'����P�6�"z�6���?����aF#3��|8��?N�~{��;6��K���14��p��% ���8[r��N�Ȧ�B/��W)���e��ckm����"6I��ߺhwFDD�WEB��(qM$2)�X��E�/��$j?0T:9�TU��0�||��M��sC����(e����jZxU׷Q�
�}��i����D�۩a�� p��	�SvG�'<��ƾ�ãV����	MM︤е��Xp>��%G���*ӕo�"]�b���Õ�P��el�{Ԙ�� @2}�HI�X֦����ݱ11~7�;w�����YR���q�����&�����hn��,��Fg�؇V�S�^���>��.���4�榤}��������Ot�"+~j����"�%�`����W�
}m�?eT���u͝�_�Z&L�F��CDL�����9A*pkkˏq�pq�⡮���?�xW�I�v�SR�S:���J R�U��0�-�u�T��!c\�W@;Gj�p�Ic�tdd^��6��H?�v���_c����Q�C�� _��\mh�,,ts=��D=�T��_��+���_+��1��"�.5Vѩ�0�9�HW�
������NŰiL]��㝳��ԓ߆T�b-N4�X�!�ѥ�*7 N8h��׹��:���0�OOˤ�_EtَD�b��ţ|b'�
ޞ���QȐc�7�bq�b2_Ǡ1Nhc�1Kp�,�P�Ģ���o���F��� R��r�eU���mWa���Ƨ"�9��+k��uZ$�*6�Ud��Y�̪�a���W��b���K���t�<iק�)Y2�p����Z{[l���;=R�Kţ;|6��x�Â>��&�h��L]Q��ȒQ��W��\�E�����8>�A�����,`�E�� �y��7����YQ,�˧6&~qk/^���m�(�M�X��O������_�.s�E��L�n��PBv�l#����c��J�&�<������,������>ߧY%t���T�>�K������&t9
��چnA;���	����"����?]p+��hm!]��r�?_I@9u��g
G��\#��Z:O��0����5V?_|H��
v�x�&j�\ϥ�W~��s���z�ֻ�!����	Ve[�Su��梦���{����z��l���kr�V���s:����G�M,�<t����ю�a<`%
�g8�/�lG���'���n��.���y�y�0@�Ȇ|A��[���_cbR��"�pj�;�=iD��YN�Uv�����a|?<��1�+���ĥCA-�c�ig������D�DDV1�-���DMArѿ�_�m*���������²1X�M����X�t_����05��0~Ã��<��m�=;�M|�1y���ъ��݇fB���f�R%�Ye��4�i�S#�I�{�y��{���ȗw�#3U��~�#&���ԉ�ls�S�����Jb!v�Ϋڨd�{|��a��b<���0
��o���ajb������n��
K��gr8_f��/<��W|���V��20�"O5�T!6i[m��Yk|�Jhy���H!x�%�A1|*�v�C���h�h|j޿U>��Z���'��[��v+�bnv��@S����Q.J|<Mn�";�o��Y�|�[�o�h&ȩU��Tc�p,p�Z��ҼS9|�B�e�:=S�e�o^|�Or:;;v��I^��K�5^����.�͐�ު`�p����E>�á	E^�a���0~7�A}�e5�����.��\�dHu�3����ol��b����1tl��I��?��ҿc�ś�BQ�1(����"Y(��W�����=�z���7�Y��mN_5{�z�,
&�������9�\��і���-1$�ez�M�o���E��{�֎Kߞ��b��s$�J4�v�?=ɀ�N�:���Ԋh�J����Ս>N)�CJ�FW�%���iq�t�0/Z����0��X_b�ǂ��4����S��J(DG1ĭz��.-��ѧk�qpK(1Q����q�]X	�"�C��vf���*�Dy�`�����ǳ�!�-ň���C�/oq`��Ia��f�K��4�s�:�^7a:"���\�+{g���j�G�3z��A��+?������h��M(C��v��[�NP-&���{�e��O���q�!�9���>��>4�WX	*I7�;��݆���V�5��� H�*N��zB�I��}�Z��*�n�ӣ^fk��22�;�iqf���O�n�%����$B_&��W�������V>���o�Ҡb�W�&Xߙ6+I�RM(w�(A�`'}7���t+�sC;���x�������.S7R����eQ��f�&('�
�� J�&����FM
< ����U,|Θ�JM�_;�p;�;���N_�^T֩K�b�{AU��6�1�.5W|�����|��WX?��՗�|�N��y�lyk�V�����w���H�&��W����VS6C�+_F�}���5�ɪ>m'�Uźi��9X:(rJ)�����w?��Qu��!>T6�.�DsTr.jvt�|���k�C����\���r��~v����.�B�� �G�i�xJG��˗<3�vv�F�A�B賜a"Ga�_��ε4c��ɽ�:6�W�M�˵��B9�q������~=M�n��8�a���������[�P��
���uh�����A���g��vF��zk�/[��aM�������L�sR�ӏ�Rԯf�T0wE�3�Ԣ'�jl�;�0ˊ�=�6�3AuH��������0�7��F���XKX|E9#).'��FK��
װ}S���nǂ��,��jo`�Q��l+*�f�N��ox��x<U�����Y'��2�P��sɄ*��]SַHf�t_�!ى"B+ђ� t*� ����W������7p�_K�UU��Ⱦ;
�<MWZ�1�r�'���$��R�E����1D�C=�Yi1����U���_nC���	�d޲��?�h���:6�QJ8�vB`Y�CjP'8�̋���%�D<��2	������:V�`��<�#�<��P<uK!�$�Ԍ-��ѫ��@>@�v:��Z��n���a�̆ONl�_|��Ϭe�2��BX2Spn	z8H�P:��r��N@C/V;�R��9-S���|�W����*	�m���
��9���!�^<E��#9�%�!�qn�Ÿ6&�4zU]7K�yQ0��ͱ��?n}^�WW3O,�K���7&"�S�#�>�«���p6�LN���/�2Ďywtq���$x���S�������zh���@�ʾ��Ef�S�Wt��z�e�A䳴h��F��*���a�)(��
�
�mT&��M�o왧8������n�Aɍ8{M�6�Y[�u�Oq�ᵃ�A�׌�ڴ��RMK�-I��m���ϘõdT[��SW����t���*N�-�ҋϲ;��%	ג741[�y��h�"N�,�_P󣄗�V`:��hS�xQ����j�k9��3bCHԓ�{Oi��#{��dm�O��	N�<�m59զb��#"����ܵ�q�[g�x>�M66��ZC�h6��?]�K�X��c��ta�p4{Le1e�i3�<�~�8{���g�,
"H��Z-[��+*�3\��1���~/�s��K��Z�#qܢ��&�����~����,tO��
�0cبu/�(�U9��Y����Z8���һGBԭ�g�v`��$M 	/Ơ�2�K������N�ևr�ބ�1�ī�,�k6��g�^������c��%x�//EX�{!h��t����;
01��,P�<����.p/|� g�t��q�)���od��em_Y�'�3l?�熍���4�pm&cĘ!N��3G�ێ�����s�j�3�47���~�B`Ts�b,ω��-����s|l-��r���X�غ7:�G!#��n.y�8���)wSj��C�_�*{�1Jʟ��Nn83�sԼzы�ɕ��F��Z^���K��Q}�i�[  �l�$/m��D)�HH�YZ8�}��]~3�=�"
=@�q�����L2e��PF&�cr9q<ҋ��d���-T���O�����)Y��0a�g�ܟs}ρj��`�!&�mX~��u}s�"�M��n��#ꀺ*���}y������s��I�>%J���d�_#�=�a%oV5������>�P(�ph�˙?��K�rVm�/�Q�g�2?�e��gɏ
���xk��f�N~]�����hE��2*:XF))9#��p���bz�3�|�~Z����16���`uLL�_�����}��H��^���L�}��/�!Oo�?�Z���n�����kG�_qW�}�V|��y^]���t��Q֍A ��領>{I�P�c�&�"r��,�R�S�{�=^��?^��q��[fy?���k\���r�|��F�]�ߘ֤S�_z�6�h��5���S�v�qYzM��o�5��}k�noǙ���Y<�C�ƕ����/;�r�T���Զ������\9�9����}nH9^y�O{=à�'e G��|s�iɴ����M��f�_�X���a��m����r!.d��C£a�[x�Pռn���[�b<���L{���Oq�U�:��Lz��F�U�9�$�:�m��#��M���Q���޸Oدm��>n���[j��Q����k�f���6cbZ9�}CU�:�s�vpJ ������s���oƄ+=y���W�%Za��<Z��ڹ�/2Ƒ�K=�^�������gJ�V���A��v�����K�#�ߦP�Pf���p#U��.2�ϛ%n�TsNy�v��~ͯ�w��=�f[�p�<���>S�١s�|	I�&ˡ�P�	�[�\u$5��1߫�;5�������}��;�l� ���S�jGؙEzI���F��2M��s�7�9�/�d�BBr"bƞD�A�Tn�V� �}��t����s�)�
r���K���F�����H��hDov$ټ�,]l��>�9�+۠����z}�n�H�ȋ
��ʈ-j�"���qAl'��%gA0�ϸ���_���K�tt�_;K�*ѣ0�dh�2X�ęs�n#܉|/7�@ =
��
&��G�t^��:������Pa.&s�:F%!]�m;��pc�[G�'&�\�`���J�B�X[ִ�7ϲ�^�H��+}l��U���;\��rg�w2��[<�b�;jo���=ryCg�-���d;�q����)�|V-8hޥ�C�,�XVXH�zG��I�.k�4��{��Cw��IG�篫qK$�RT���oȴ��%X�u�2�BE�#!R���k�J\{@��p�	����(��j�9�|���G����Ifz���V�곾��ϒ:�Z5��n���V�܏]�ֵ�_�a�����lN�f+�d)�����(�o����C�;��Ȭ�0���k�	��_:&�lcH��ly��:�~Cn0�޶H
���\L ǁ���b( vlG-�w��,�������_�<�����m2�;���}�#C�v?���9�K;6od�mH"ÅV_	[��A�|��l��'iD|&mn>S��j޺�����A@��M-ox��v2��߭0���v	���� Z�՜7�dnP�7�|r\
e���f�F���I�>�Ev"Z�$�e��9�O�8^[c@0��0�UU�l򎸟�"����������酕ge�/�Xj�q�N����X=;#�����rP9s��=
��~F�U���q�dd��Ё��o�����v����ԠayRjU�[X,Q�D@�O�Bd�=��l�fF��u#�� 6O)��%���_c+4�-�E>qڋm�������8� <Hd�߼ϕ�Q."q� P�s�pG�	�#̇�wq�x,�Oi0Ϻ��7Bf|ۺ����*Z��+�eQU�";[�=���f;�3���-< �E���p����( Ԋ�E��J�]����ec]�B&�++6D�d@n�p�ĄH�V/����9`m��˕�F������hkk�벽@���<�
ݢ���aT�0.a~���V�"����E��iPnp	�ǭ��beU��+���ddH/��I���?K��N⯢I����DU�eR,*���8(�H�j�

&���~�c���՜��7s-^,3[��6[s7�h�,h�5J�9��
���k�*N�����3�P��)��C��`�nYD������w�CZG��jk3�j�������{Wb�4��`I����B�Vz��i�����5����G�D�t1J���$�f�5w���M|v08:|�����t�7��p�A�R'�h�d�B���(AG	����-��-\�FA�b��j@BԵ	
4�˝�V"x`kB��]��>)��;A���0��A߶DZ��t�@C@i�C�_�*��mmS離��i*��-���qI��NS��Qx�����>�TIB4EC%q
��=r]>&j��Oh<�u)c3V�lb5�S4#:~Q���}�F%���R��u�DQfG�Ǻ�B�<�c��	�1��^|�r�v�X��w�3*��V�����BPN��<fY��=d���U���S�1��t�K��� �Q�l��J����h-%�CWH�~!�*n��v̞��ݶ���MP�ٓ���h�i��]�����Mg�ITÈ1#XX|v���j��lE�r���,L�Y����6���v�g�������D��bK���J\�M3���q�H�~a��Rx߾$�3Z��Pm�slӂ�O x��G#����u���A�L�����F �C 0�*����� �]�.ߋ���E�E�:]e���R���y{�2��Όߓ��x._�z�At�f�|������'��!��/�%4<����-S��A%��冽y�R@�d�rL��5��E��BlR`	�|��5R�^�7��l�1�w)Ӡb}�0���GD�}ng �Ɣnӧi�F�l��H<��j�R d��$R0�?)t�1�=O���7^�╍�2k"��џ<�L�ݿ�Mk.o\�Y[.��jY*������a�M�M2ׅ�$�~!�	���0�Gy����]�br%/�|��^;��(�� &^�<��1��p����Z4�`��F6�T7�k��G#��p"�D QFz��j[�z7�G��n�cpS\� ����&^� ���aM��k�D��v*V�@�mù�("	k���BS���od���q_?��9획����OP�B�I��+rY�(�l�:�����zL�"O3�*����qZ|��u�/f=��`�b��@æ� #q�]k�?a�)~�򶱄�h0j՝gǮ�#vIdShIs,���˗����A�PDz$�~�%�����p�-�C��G�����w~Hbn"+G"$�w���_k ��[d˻�����a`l�����_!�����Gf~0�/g��[���	AT(�jú�(�U�l��g4��ul���+��^y]֑ex5��nLpǐ \"�.���u�RYLA�, T�3.݆��Z�q5(F>(���:�|@��ٵ��}��[���LN���
�g���	hh�ҳ��t(�T�HI�)9Wq�����ק��IP����V��ܡ!!���!:,�1�	�B�zj6�^ ��c���I4��x��$�4���O�k��JG���@ރ���>�K���ӈʅ��B;u��{
/����S2���B/���{��	_n���}�����
�d�T��ٳ��?4�@a���]��*�(������O���T�ȑ��`�HU\=yr��Z�X��an��CdD΂�����4��5�#J�5C����D�48I�]r�n��r�x,�
u �4�w4x��"�X��S��*m4W8- ��$��+����}^�.}���"��l��S�M��pP�N���H��+�B�VbKq��������Ҕ������n�.��R�b��V2@G��=~�a �\-�BA���b0��>��� 1���5����A�����sC1��� �D�;�7_ r?m�4��~����7H}fx
���~��Z���~M��9��.�*�nk�x �5;�&�y��*����+�`�T����K.��oD��x�7$�ut`==á�b��R����t6P��Ǐ�B����q��]��'_k�R^����1Mz��z��Qf)��E"����4��C0C�>�<��yE!���rK`Y*�=�$^����T6�Xɗ;�%�JA[Ԩ�[mH�m��Ph"�-�$ݗ<�pt�)H=)=:�d𨎿N
1��߯ 0�Ej��\�팷q�q����s��p��.�~�b�y`Aa[4�J������"Te�CP�����"�9~���=��g��9Y��B��[&��Π����e�o�����-�3���ǳǾ�h�UE���9�
�ʐis�Z)�#�-h�W�� '��]2D���&���Gƪ %�02sr$��(i�d\�
�1ެ5����(���X���ڟ$���T�li���X
�R ��"�o�l�FrPQ��m>\�MW����l�cn��e6YT����_I��8�����ⴊ�:���)t�tj��"2�J�ۗ�ǃ���������Hl�K+~@΃�Wh}�Wa�<�4 ۿ�ݲ�3i�"�C'*�DT�^i.ܱvۯ���>�0�B ���z����=��:C嗣&�&>��C$iy��>�<#;x�vwե����@�]x��#���<孷���j�x������f� zX�S�aB�&u �z�!�V*�$ UO��b�X�Vf/�l���%�alBF����騜U��gi���>4�kjj��Q~92�ߒ���HT2�e�.�X����# J�s��y�l@�4�. ��4k�&��>hd:� ��6H��e����h&��c�T��b�9��t;#{���#��y^J$n�h���z����J�uȍ_ݠL[k5�e��qH&zn/����A�|�����������<��a>�ջ�l�f�}��py�.l���R���j����_8XW>!?��$��i����s�)Զ�u�+o����6 N	�s���ɀNl����l�jP�K3��Zt�TPnj��g��9G덊@e�(x��[2-�HY�9�Q:�I瘠��:1ǫ]�G��0T1�T�z+��zf�鿻�4��٫8��K�~`�F
F/�0!"g��D�����}�5��Kr���3X��	�2��uv�趆��S9��A��Q��Ȅb�L'l�d���~�]Ҽ�t3�~��O���.�>H���>9�Z�j���l���c��l���؛zq3�O����f��o�cي(+�~��gVB��2�K�)\d~�HHA���|�T�%^
0g`G�Ĵ�C,��B����[d��e��w����w��7���1mh�2��f(���Y��m��xs$����9�lr2��-��!f�!7 l��I����N
D�ٽl�7�K�Φ������oV��� �<�.�*@0�{��i�E�����\K�meߗJ����]��.	������?RPHHIHII�ʯu=D�XMՇ��ݑ���A;a��!�ZG����%Wi*�;/l_֐R԰7 *$OE1O�A� 3�&@M�
{�G4sds�]�a�VE���
������l��� �>�Oh��eyPJ]��]��Q[]�,��o��b��v��<:e�-W�Fɚ]��[�a�Ҹ9[� ֪�=��Oz4#�l�lRX0�K�1� ��z,�4ğr� h�V��� ۏ�"�-��v7)�Y��zRH>`+~�wfO��A��#*_|�7��wbc�I%�"�h^`5Qv�{�б�����8�e}����׸#h�/:����t냆�ҲI(p���k'�&�^-���H��<��}o'��S�t˟tuu-I�ɽ�ɋ�P��@��v<C�b���8�j��d���ː���w�j�4��ٿ�L�I���m0$;W/�1�@
A�V�p>2<,��H+<-�Gl��hM�'�f�)��b��N���#4m���8����B|���K&��t�8�"� 9�L}� =�i����+�b4���\*߫�]̙;������h�ɐic� f���\H���0~#���:��[Da�9�hSq(�Ua1��R����1����M}��@�5g�&� ��m���'<���rn���oR�#��6RZ�룠9�!Sex�p�C�[hwh��UX85'&���'?�����$���:x��vҐ݆�mG��o�H�|E���"��X��~��l�``�@S�����h�X��΀K�$Z��s�X@���U�H��br�����E0/!H �`h�3���a�ێ��O�j(�P��%6O��IE����J�� �0�p�n��u&�Ā���*�}
H��_ł+!�m��݀��*�c�@�+�7�����l��X6˭<�;M��$�n;�e�x�Z��g���ԧ��Il�+�F�m]rh�� 4C@AF����a��6~8
�#`f@�7�)\0���4���<�P �$��X狈^��a��� ;��n�"�l���-�yy��G�dn��� �-)�~�r�x� ^��?ˬ�a�i ��Ѐ���L�138����4�����j�Ρy�l�h^��������	�J��6��Hb��!���`F��i����W�7E(��Rm>��� ���^d9�p(wt䙙~�LGճ�d���	A��ܮ�꽏�����{�;mp�6l�R�1���2��_{e�Jv���(���{ ,�U���!����)�X!��ܚ�(;�~�2!
�����Iyq�E��ݍX�A���C�sw��\T�d����~���9����5�)�l`��90����כMX��[���r����"�#ض̆��r{:����^��z8��Z]�r>��|�
���J��z���ɝ�H���������_�X�x�p���>V�3q�S�WP�T��S�����v����L��f���wu.��V�{�v� a��������g�L���gVi{��,�X����9]K1v�����κ��l,���:��.ju��d��&�Ϟ,2���]!���i�.R�U�i�B;�mFf`�+񽮸ѝ�u��q���Fh�c1N�n�Ϲ|;?���b�i�n}�	���,c����<��O�$��|�5�ި:86. K��I\Q6�yc	��o�r�(hIƅ��A���W�����}}�㥠=.���������m�M�
?���;?^��U�G�~QR�����Ix��	�[���+�_c���8!p�9����y_����cp�j}��p�PU��if������4}�������y\-X~���Q���@�ɝ���+���_j-���#�.R�о�[mkݶ���P����G߉cU�dBǎ�����t~*�_ʨ����o9��M�� �g��r�w���5S�xd�M�����C�zǫ�A��k[��w�H�Fļ�h�Iv2�^�U�+�Ľ����^��00���k�׉)z�F�UI��F�=Ӷ�׍hw�=���\��5dw�v����Q,���r�����;)���� ���2���i[�E{�|;�5^�����9�)�U�-��}&ZS��k�z��樿U^�~�dp�d�r4��u{CJĞ���v��nG����K�����:���@�s�{G7�:���v����ކTW[+�����Qu�[t�I�jG�s>�X�ٮ��8�hEn�~�pGl}Y�_�T<�{�~��\{Y�N�&{�� ����dx���Hq|��w�_�mџW�OZ��%�=y/%�;����W]t:���ӕR�ΰL|�'��P���r#�-F����5u��7Ew{A����˖�� ��yΆ蔲�k�b��}�xû�����Ҏ)��\s�q������ֻ�ޮ}7������:��'Qt�V�7�9WB�O��W��s�.��Km4j����lfD=�MR�6j_��16�-���[�v��7�ٵ&>1U.{��T��AY��u��ߛ�%�h3j+�������'%2��:��X����kk�����KB�2�}s�f���������'k셣k�4q?�8���J�l�%����*4���6��aN���6�P��<wĮ�� *����*7`��$,u~�p�&��=���B��/�;"}򑢵����*=�{�|ԅg#�Ѱ��-���%�$�H<ߓ9!�fd߳.ץ�Y�fd�W�$s{J��AM&	pG>>4W��p��k�DG�l"nsE�8����f�M���3È�' ::����!�zafn!p U.�������f
�=, �+y�e*zW�g zqc4`!O�Gs{��67G����z�&-��r^J���+�$ex݃� 6�_��;�|�}|��wW5p���?�;��+\Q�h��K��L�N�|��滸�5��`!�޾ߴ���d����l�8�V�{����W,�]]��u�����(*	Z�o��NQ�9�/�g��6S�ÌA ;�fM��3$`W��\=XhQ1B��m{�=�:���$z_\i�{k�E-�N�ɣ�����,��:������L����*��E��;׾Q	�� ��(�8(�G<RXI-�S��ߒ�6����4�\��j��|����CL%1�,i��J�sP7	����>�i���R��K����ۻ�M�)�g��p�ܟ$����~�/���z�Fݥ��HV�Cj1@
�]d����V�W�I��l�X�
)�np��\�l�˩��oT�aaV�����	9���Ȣ�~����`9�Ǧ#�M�Ǯ��.BYu����������cH^ �74�g ��eEFwzb��7\R������W �$-��κ�D L���%b��	5���n�&�[Z;)�$1 	��3A".�[?��
s�^;��/�Y�@x�VR�����0;��/CO����1R��
�Sw��8|U?�b��g�O�-!n�p����灒£�?����5��fx��4y�g�Z~��yU��`n���=��x�>��¦�*5M_6�﷿�o�uO8u��OuE5樜>b�94���+�n8c���+R{��|�V~N��j	9~�on��ڃ���ѝ��Jg��(�%����]U��yGc�[9`s^nJ���'	Ԝ��6�t8�Z�ޓN{��6����,*~
�̸�zƛ���P�H.`Dt�vBD��^��DI���S���-O��PVڽ`k���Y��C��Ư#��w��ʮ�u�,�P�jGy��ߏ}��ke�O~�捎�6�5�)�֢����zG���֚�����B�r�"XQ�o��uɅ1fXo��PX]�[��7l��pY��6�I��w�i�z������v��J�%婻oa�E�=]�.�~�G�r�?zJ��4r�H���i�00N���#�,Q#·^n2����6���8 �$B�@�L�}�b�^W��(��}~��dZ���s��Ni"��Od��I����%�8���/O��/糿���?�sK�~w/a�e6��U.�"
���n�ϒ�hh�b�a??�\���h�Q,zG�S��`j���)�~��
Z�y��fѺ+����#ꆸ5�ݤ"������sLWy�������qP'3�T�F䥝����(�4��X�~��l���ğ��t�,�V������]�����W��G�85M�.�F⟠�heU��p��}WUK�?�ե������P�U_[ˌ�v���.b�+n)�n��<�]��?I��$�@�V����uճ�(�?~7��L��uX<�p��7�N3k15Wk�[��Ѿ�k��j}��Z;n�h�?�н��8�e#���+*ԏ���Y��/��N,ե��ȼՈKm�G2KҎ��������3Α��?��SRo x�j&��Y�������1�����\9I������Z����:LPЂ���"�>U���	�*�����O���'�ӛe�y��}�Km���gEX<H�w<n�8c4�eE�H��������M���XZ^�֖���=�3��P�� |��������NI����ZoT�G]��kn�6�t�ܑ�Y�����g7=��^!�늀T��Oq�s�B����$��l��c���/����,R���ѼՓ�]����>��3��(�[a��@܎�/����N	�3�}� -^�h�x~�� �Q	��X�%�/)�D���ao��S����o�y+`p����8��Z�΄]�ُ�؀�:�%���6�.@S7��G��H��.Ȍ���<@�J��e�A�>h�#�'�7�;�ǫ~�<���+Ϭ
_\W�~ݬ����'�~ʓ���l� @dx�uk莑�9=�]�v=sH�����m�ĺ�%�\����4w�Oy����g]xz��48��`�[�nI9��z
,��׮�]{�h��l����o���v�����޿�~�ޘ>�^�Mx��i����W%��ȍ~����p��)���%Ĩda�'rh10-M:6i�� cfA�)%5���>� �y _/ ބ��N�o�1�r�dg�o�|V��5"�ܗ��]�k$y�2Y�Ji>�#��A�.6�H���_�]ND�H�~&����@���@X�����T���c6��fܴ�R����\�)�C�l����z�=��QT�\��V_�x�죵����i�\��.�,�f�ڽ���2��"0����&�Um����T�OdL�S��dmMU�Q19��(�c Y�<����<��p��w;��C������bzV����|6z��Z�0H�AW!E,�8O��Q�F����Qƪ�&,P9��9ƠkA5���rG���W�f�r��y�jp*��~�%��CLP��A����|w�����^��+d�C�~�	?%��d���+e�2�I�����o'VL�U�M��W�?��d�]�{�1K�i��J�~8��sᚳ��s����N����h��{�ㇵ�������{�QA%DDZAJ��K��E��`�!DA��`讁�������{b�O�/��Ď{_�u_�ޏ�E�WD��Rx#v�n~�w�I��)��tR�m�}��xFj�tߴz���,�%.�[�@1>�.4~�-��]�g�uY�d��؁���|BYfB��?�,G��{Kf��d��IG6���(g}����"Sީ�t��eyGz��]]�^�~.[AAM�I)g��@k@zԥD�MQ��L��b���c�D�`_w6�U�f�����9�޹�ܪuW�}���4S�"�L#��J�#!Y���r��;>O:���E�%=��i.k���=m�@�1�ː��:46T�@sQNoma�^�M֔��i=�a,��;h�AY�8��M��@��pM�������C@R�j�>qZ�j�$�i�����<h���1x��L�pM�/���?��K�(�^^��T��r~18��~� ��#�HƵm+��F�: #ؑ��0Q�6�P��)���W)&l�_MT��,�0!`kG��^�������w�����i:��,Y�]���D�(�m���I1f�K���|!��"�e��ȝ�	'�WǵU
�r�ɶCЧ�z����@2d�3���BuV�n�}.����]�1T���8Ʃ&k�>���Ī0I���ًY�l���9���wQ�K˔=��-�x[0�6��#w�����KX���_T�f�S���i��#����_�x���(������O�~e���<������7!S�xSd���B]���B�l;/[A�;oWۨ�t��ݢ�����[ߚ7���9>��24$���G��O=��D"�Yyޛ�2kui��b�׶c��?��Iې��yr&��&uT</ ��"�o����7�}.'�j_W;��H�1ez�E�)fd�E��	�͋�)~@'�ǫ���z�Nļ�!j<��"�@�����۩Ǜ�i<[��_�}�J渗��-+��g�"�Q�vIVWF������C����a����W̢�Z�|�&#�p���X���rb�˚�=Å���e�	��'�Q,L;�[�2�_uE>,����}�=�Lg
6yx$��4�$�5k�A�8�|���]����&�,]�c�u�w>����.�~�ъzM��bi¹[��R���d|×'��(ݽ=��䡯�b�����7N�)~�I�$_<�rW�u��划ĸ8��Tt/w%^��N���A��bs�?}�"�	x`�ř ȍ�W�����&yDh�_��:n�����?����2�`��Rx���-G�S�Ǩ�L@�Ȅ��i���p���S��@��j��Fz���Ț�r�P��;��|�w6ў�r�NxkBN<�Z�NtP���$�jvH>�����~���`<!���ne���ځ����@�����]�:!B�1����!�s�m�Y���r���È���mZ�Z_�p}t�ޛ�f���9��"�Ғ\:�$O��pg�>v����k9/��B���E�k��Ne ��(�`v�E�$wt��f^�]=U�Ć�Q�S��g��F�ٳ�y0��ލ���h��1n�
��N��(E���<��7~$����b���g_O/f�N]q�hH[���M̆�# ���� Ͽ���]��>/���%����EAF_����)e&wa]hI|h��eߛ���gKk�J�mׅ'������ќ�%�PO1��g�@��2�J<m?��F�7��t��I0���kLdr�~U)`s�E� Ѩ�{���jIɉ=edXʓ��.��jq�����Ͽ���xH4�ڨ�1��p�V7FO%\�!�E�̑�1r�3`4/h2��������Um��)�R���ߢM�_�}�S��Ҿ��kbN��[�T�>�-/z����ђ'j��x�Axη_��Ʋ��a�a���^V㔳f$�h`��׍�����q%��jT�L�J[d�t|���*�z6'�db�/(�'���d�d���7�`:q�e�R7޽[�ʲ����Ҧ'��N��#m5"9���0���ߠ�\��KzG���G�Q���F��b��Bun��Rq�J��s1'��3z�(8b2���R�`oX��q��
ὴ�k��Ϳ��?o�a��\�3ct�a��Ez�/�P�(4���5�S�7������]�>�V�T�+�Da*腡��̊=N(��&��8<H���Mdޅk)�n�l|{�������{~�����[���y�X>Y%�����Ԉܯ)�I�\'I<�Cwv♩��BN�����b�ĥ�]A��#Rb�6���[0��n^�
��r���@�)tnӛg?�H�{{��I��/ͺ�`T~�ۖ
\ڮ�-W�|r��,핿c�X�哗~!���nS���ܼ+ho6da^���4�#��n~O����K#���`4%��溧�8�Tm��A7փ*�5yFV
[����Y	i�ya>�ˏ�4]A�������Hp��i0�YE�{��,4�ڗHf����LÈ��;,�� �J}+OQn>�gh��xL��X=���{j�+#��ry�]gՎ�rO���f��BF�|Ԍ4��H�li�e���%�;7�cr*��疝I�W�or&�8A���+Ku$;��7�RO�ao��lr�!	�|�d5�몮]y�ѫ��d�C.���;N�'w��l&�v_��{�K��f�S���/����WI��X�r?!=dM���X�i�.�����I^�.Hg�X�9��rY�+�S��T��g��L�wc��EX�MRV:������lr,�.��M���3N��W��t���T劷�/߾Q`
"�%%��S�u|���{b+���/�dz�6ș����ʓ�
�e�T4�J60ٶ�$0F�#Ll�C�\��^a�,1�'tҖ���Reu��mn��mޟz�M��od�7)�klu�~��_�X��4/�������p�D��u\_z���I�W��DX��HWl��rto�o~e�)�lh�96�$?��F�^@����م8/;�ћ��\�k��r�<�m\f�y���'C�*5;�:��7I)����
qtY^�v�X���<�� 'B�1�V��w�{s�e+�x��+��TK֣�v�e��r,<=�$$$�#�C3W��m����^�����J��UD&}��������Ok񬎑����+�!�dU��Zbo3��������U�Ӡ.�@Tп���?��n�������?Y�n�w�i	��pI�q*uv�*��	�l
M.z�"U,l��c�l�}d���6	Q�#QHv6q��.��Y�daN/]%\�k�F���[��:�$�K�����Fn��Yh�b�F&���.�"޽,q��#DOm7�k)���6��Q+�L�(#��(�Hg\y��VE�H�S��'�?ޫ{Sȁ�I�S�F�n/N
��&�Cf�ɷr�]��a�_,U"�^��Z=��r>�<+z%xr�X�5�0&Ȳ�����p_`��.(��o���
���â?��2D������7�V�/�����_�ܸ)o3k�n0�>���W�8�qB�Ιd� ۆz
��	���[o�T�UK�o,��ׇ�v�������W�,eb���W
9X��%�b�aϞ^�"�(�!/}�c��&��M�7.��|n5�?�F-�E;�b\_�*�蚳�5.���p�=�2ȎR�ݝ������z� zk1-�y?�+�E��a}
EC�M�'�n�+^��3����h��hA��ُ���>6#[UR6�9J��D)�19�<&�kC�� ��ti~m�u
��X>�]:�mۏ*��_$6S�9��?���=�k��N�+~���o���*�53W�ޫ8v��L�P�с@,�����h��jج����
`dq��8:�s;�=D/$的<�*�����JTW�y�V�* �-��1�H��29��M��(@;���� ��4]���7��w;v�,	�9��}��p�*<���p���˛K���89�����u���7��I'_Zjn����ʖ��������$+{h����tBI|Lx�ى�r�W���˔�P��$?!]=���MY�F:泰�2�>� ��Du�M�tb�rr�VnKW��S���,ƕlUفD�GS�;۸�&���������5�5�h[H�^Q���O�fMO�-J-(J�ƽ��P@ (p����ξu�V��~5c��/�ˬ���f����v�*w�ᬩS��=���}���?Y�q	��U֗Wg45�P%�Z����]�p?�����Z�~	���i�y#����(�~�y��K��^ڮ,HB��H�9�|?滹���s~W=�m�$����i��Q�]^5z�c��V�'���r�p�^v�5�z������>��)��|��(o'�wR{�o��8��IИ��I�r���ξG����u��ۼ�4�l�0�+��	��eD��=@���V#8w_��?*��_���7��ųr��0�������>�Ye��WTo��x��1��%�� �(�`�z��/sI�D�o�V`U��3N��쌉�u���5���ŹĄ�?�BJ��~���ؕњ�;2��Ns<�Z�y�i���r�_�)r�~��n2�2�SC6�$җ�b�����t������(�ו��0(y�k����덶Z�H�
��'�K~(!��]��-�h�(�I|<�㓟��H�$���{y��j�����-CȄp���[���Ȃ��"�>����SX�\�����N*Q�ȴ����b���[؞�����]c;��I@O�����0�̭�K���Z��&rٍ|�JXc�L���-�<��t���L��������8Zۤ0�y�~��"�Ef�ۼ�xc��r��<�̬�ץ���q-�(��\nc���d��I͟z�4 �8C��篸tH��/�AP>�ii��0�I�SWEw�������j���(	M|��+���})Mr�\\�\q�}��ȝ���d:�{h�V�.�h�cx�#\��b#����|�+zCB�[+Ȼ�>���W�G�u�LT��)��_A��@�|es�n/�cut�:'|���Ǎɺ8�~@���zP�j��ρ����׼�O�b�R�c�����Y����	�o%<{�|&Mwo�B��|�g.d���(6 �9��i�!h;e��KbM�������"�ک>-?����t���Y-�=QQ�4����iN��7�(b P�s��ݺ�����fe٪��h����H��Q��ǎo5�6��^�&�)�� �e*��.���6��OҨ]���0��#b\� �1���*�?̂�1�oS��ϫ�?RB:�.�k��yR��[�s����=��7ys��rj�L<풐6u����zn�>)�SlQ���_�[:����uq����������_�,���eH�TB���.!|3~�������e�SB<h�`?��*X�7��3xD~;{�<�M��M�0�4����/ �qdޟ�ؕ��W:�'��ZIAϙ���hh�����2�"?n/�!#�������Ȅ���>�ގ =�- X�է#u��_EJ���c^�r��wA�	�$ê�>��J2�.)��L������`����l8].�֪��[���7��W�����k!1��v�u���X�=�{_'�X�뷓-C��N����g��
�U6?!�Z��3x�&)��^'�����xFv :�/E]��_k�\�������S��>�9aF`2�Q&i���_�-�o��mR1KS�5Сٝ�	�|����lO����r��Xu���>j;}�����G���tBE��	�hzP�7�@�i����]I�]K��F��̭9�W7��]��3h����}��mKww����SE���Q�w�/ۉqv�\K�b8��è�52��=� �|������Ƹn�w/���hD���	��x	}w$��MG�vko�Ę2m��7L�t���ӿ�Lս;�t�RK�&Å�t	�I_�ʹ�V�i
��������V��x�x�jR�f!��~��C���̇�q��0'�������a+ϳ��})p/���U@
ܽ���<�
b{ �V��-ZB'Y!�w8�v���A"�p�T� �D�w5�+D��g�[��۽�Phཅ`u�Ut���T�'ٯ���- $�K�7)���8B?HĦTﺎ+�
����7��Ueܭ�?$���p���~��r[�W7+m����`�ω���@��4��;�ܚ��8�1�ʅ"��v��^.�/1YAA:�6��|:���

�~������Ns�S��gϺ#`"%�/�� E��r"�v&^��?~�c�_8��,�J�>%��.�q�����Ϝ��]�� Y�-7��^���Zz.WZzl	��ȱ�\�b��è�uC���s&�6�� ��=|�R������@���
r0�lu��IF�?=fb�R�� � WzH��JV:7�E��q�W�&�Rv"v;��;�3����Y^��<�.��(��@�䂇�F]�J����f�?@w��(N���k��2r�_�� +��,�С.�q~о~���V���fN�6�����NG�'ci����VR-`㸫���te�Wg"upɣ��Ke7�ؽ�q"W�,p����ʽ����b}�k�H� ��C����\�����wo�Qf+4��"�-���K;5��tq���c�J�|�l�Q���Y����t*I-H���zO�l+K��h�UB�c���ճg���\<�r�rS��}�H��n	n�U��~����b.g.��je�B�F2b�?��%�n�\�tV��UZ�@tP�Rr�ټ�!1 !b&r���Aů�>;�ܘO=�'�_<��p1�������ݐ!;ܪ�vn��80h�q�m7�����>��!lW��kUk�<̣�b,/v���`��S[�:G+��P���F'w��c <Z.X�f6�`1!wْ��Td�;��O۠}Wp�EC�~U��ݲ��UE��z��7��/�?M�M��El���C����e�� �� �|8��!f\��ʇ�J��aѷ+?����M� ���1U��EXCsপ�����;�e�Q&)}��m>�w>2�q�����C_�P-�5Ir�]�o�I��[�!���!y�ڵ=_iқÛ��w�Ol�VI\��[���&��C]Z�;��=������^С,�à*A��>`�?
����Ʈֱo��^�+�.D]L��ȔM��C�*@���G+�즶�ǒ_�.�O��{}���u)������Y{��(j�c?���u���c�����S1���^���W�ٞC�ղJ"^�6����[�����J�2��z)}`�j�y`a��4!�ck�6�b�]�x�"+{-A��zNr�"�\`2�}u����Z���t�\��k����i������2\����֏.��	�����r���������|��}�b��8xl}��u�
YNԪ��_B7�(<�-��;�^Oc��^�������O!��<uD�C������8��hB�``�R?�Ҭ(@���q�}MHh}�W�δ/띜o�u�U�+I#�� ��>rR#'��#G?q��<G���Kt�ޖգ��8U�����&��^.�C7����H�PT�*����7m�M��X�a��x{�����w��o�IFHl��t;���qd�]
C>-Rg�.ebe;��D�o+N-/OE�m����m�Ȃg''�3��v,��0Q�U%��6���c(lb)�5�ϬXBF	�.Wk��C�!���*A�j��č|P�]=-���^+:�NK�T�#�]�'���q{�d�L� ���VN �����>=��*pc���Dw�o��	��0o#�X��<j��(�A��B����U$0C9F'���ǝ���u�jO�N/���rYyNɑ-\����Z�d
;��V�6^דv������=!�ǝUȔRW._{��t�C�ֵ�/�z����#������Z���{�.���<M��*|��K|Z�ՊƝzI�B�<k`I`���wU�7Cu#3�%P~��@�XZ8"�M&��f:v���7�Τ�;m�������!�u������]2G�I�g���+���E�+j��t$��{*���=ۮ^����@ł`��Y��,�s�@���}�B�� .���������v�nB��5X��Ωg�9��*Gi�{�9fd�zt0[��x�`���ê������ȫ[�X����-�Rv$�Θ
�����_�H0� Y�r�_���X�D��ݻ�Ϟ���(k��Ctө��.�)V��3q�uEʢ�f��y����K�+>����]���SQaR��KQ�t�ʇˍfe)�T}u�]�r���`l�ٕ�����Ӿ��^��ʗ~���㮝a���c��z�xX�,_n�[���ss������A*]���8�x�m����7V�ը���?].�3GBbJ&'��
�MQo�Hh���8�}-�b�n�O3�ʙ
�4�>�G�̀m��g
�.��H�):=)5�c�$L�����j�tS�f�R!P���#w9U��zNlU�V��&�ʖ�/ŧN49�����E��+��;R���nE9f�����H������:�"�5�1M�x��Ѣ�6N�Pf��ߚ0�V\����p;���"ʀz���m�1����_���Y�MY-��{d�H���x2�v�n�m�4�X��s�������-W��n���9e��|�������.T�k�;�O,�[������o��k��z:�?{�m��YXR���<��K�x]�e��eɛ��s��r�u,:̮��)�'#�E��^��J�aųgTd �`�^ǻ���Z����D�y�`��sz�ۣ���g���`�V�"��Gz��ꍼ��̃
a�!����AV�Do�-�j���RPǱ��}���5ŴiJ8X�5t
E��&��t����]�R J&��eka���.���.e,r��X�2RօҴ� �E1)%�+*{�����:��0F��%r2��-	з9�7`��A���6^���f�-��p�$x���:�*�w>Yb��b��"�4J!��30{���L$GTF7\�e�JE��z}g�A,�O��L�f&Vd��s7���/����c�Ў�Ȇ0R���:�2P�y�����7�Z�&�j����
��������i��S�`_%I
xRC����hb�l����~^~N(!�\�|��ߡ1��×��A�^H�>
Q�?
�5ղ�Y����/ 3|�8�
MQj
�?�wS1Ў6��Nme�G�҅]=+�r�.}�d�CE�bQ��������0���/��S�o�񥚡�1R����?cP\"��79Tc���b)�M�k���ٳ#g`�q5�8D{�(��S���Gps(kDF��]U��C6�9�+�&+�ψ�s�k��c��0G`r�U�=D�ִD�^�n'��-\"��?5��>\��0_��N���U�ږ�ls���E��+�K�~/��Ŗ.��O!Ҟ؎snc��K/�]� ώ쿾L ��p>�Y7]�����#�q�f��O��	Ӓ�hJz�e� fW`��*�� ��,����ʟ�D_
^# ����Q�_�m�/�v]�����X�82�Q��~�f�2W�'��^@����������ޜ{u`�:.��i�z6��L��
�w�,��U��!*'��%,����]�\�{>ԋ|w�}�Bޟ�=���9. �ݝ�-Slo�+�3�^V�9B,x���x����d���5z_-K{��lt�	#J#O�ٗ�����e�~4��v9�,B�:k�IW�6����r��k�voل�*A[B^�b��R��v��e�o.����N�QV�B�,T��LF�+��u7S�QU�BnS��ߏ���nɅ4{۔
�=Tƭ+�~u*')�W���ͻ�?�m׉kb��`���+j�yŬ=���r�[���3,/y�+q����F=���T��J���3#!v��(K�m $��If�8���L�E�([J����[+S�����
��8f��޾|��-���_����a�ź�({:�(q��D��h7?)��ЬtR�9��V/�%vcZ8p���Jf�r�O�D��q���m���3���)��;�_��P�U�`鵰�u��n��l�����7�����zUTR�%�?kB&#�gݷ� $;����xX+W�ʗ�AO��//���Xߕ���p���'A��]M�	���~���q���z+���{#^��h�ī�g�����Ɂ;͗�%�� �"*�.S.kXki���Z�1��*w���-ъ鬌��P7��"�U�,p;����h�<-%
j�].4h�<�Qh��- ��SN�T0��Ȥ2csOӴ��V��_�E�z��6S�SH%�>�&�� ^h�ѻOx���ֹ�|�&O����M�`���Ų�Y���߯�w��C�}�be�w�yz�E��"atP!`L��P���Oυ=���~������c���@���R���o�Y	������r���X#�6w/n���D��pL�v��f�8n��I+�fh���9�㉦�鋯�x3we�/���~��\kR�@�<��$�|���g_�+h�ˢֆ���9�g�?�IXQ�R��������1�%������!*�t��_޴�L��}�(�l��'%X���;sBx#�ޝ�^豬�'3��T��/(\���P�K~T-��Y���y������[�X�
��]��߸إk�g�V%�����S��^1X%��W�}��<��M�"B�p�1�s���i�x�h���O0}�c1��{���b���@��Ǳ���6���E\`0d�\)mqF��#�f�������4�����ZǲИX {j��p�@���ecY*덾\�}��<�T����g���[����9aa�y\J��U���(�v�W/k�,lx0�.?�%��|Ų���gMZq����e���0�$$��2e�8"�;"�,+�-�P
������a}{��C8%nr?Z���� JKN�S}h���p0S�������������{�)B�^����HEр�ۗ*f��u_�V}@��x識	�� E3n(����Y|����nj��!l�Q1/Z�z�4~+�|l���4˓��n�qKe�(� �Vd��;��S_���iM�"���v{��=ܬx�:b�g���by�I.�X�n"_��Y��)��?�`�Ih8ǼN�?�#l��i+]�,�,�~�9=���)���b�w����N�?��K�����M��uO�L+�߇���Q�g�:)�(؏�+�>��/1m#)J�t-����iTe�˜:�eӉ����/��Aƹ5��ùF��}�Ug7Q3�z�+ݿ�}1�8�<O^��C[�w�je9��A�y<Z#I�Wr<pTe��B���i҂�ʵ�"�UӖjyZ9���yZʄ������gh1{��{aO��R<ER�c�۶�~�:�����2`+�}����]��HG�Y���ݩu���}Y}&IO��*+{�޸�UbX��x6D�V�ez��"�-�$U��u�0l���l�̛u8���)r�Zس��"j�E� �a�O-����q>�T9�w�>?��@����LL�q���%2��n?��E�FF�a�͋�[�VE@����O�'w0X��KP�0���I�1ο���G����z�I_aծ�����"��2V���g	<K�#þ���޻�|<�ỏ��}�"FV*|�]WT�V�����t=�d+A�O�i�:���$�rƪ��H�=8��h
�����teV�j��pE��fz\�Խ�n��3/0�w�J"��غW4��~�B�eӊ���f"
�����V��p��Ɛ���H�B�#�P��[��>7�����t��x��m;��ن2�ޖ� u/��KBp�)P��,��B{A��5��醑�~��ݛ�oͤ2~$�˸����W2����-��9�cRGö�����@�Zy�~����������'�Ӧd6_#3��ϗ�^o��	Y��=o[�ެ��q�;b��tQ�_��Ɖ}�+��DP���U��	���^M��PСZ2<�k[)��؅'�Y�G�1m�	�y��q*�_zu�=E�N���o���A_\P�1��3e)���=��N�^�.��r>(){~w����`k���ȮJ�YxJjWR�i.���I�f���f��'��VwYs�:ShT]c�;?W��g������������x���`����O��U"v>��`��wr�S�&r �L(��T��f)�o�}��޻5s��/,X|�Yi�(x3�+�JFfωA��S"�}�;r%�g�?]�Hq�Al�hĤ����tjv�q|�P�{�g7/�Ko�,�<e-t{��{$�y��5�����틳�%�YԎ����=mc�ޢ8�#I&�"��?K5�E}dB7<W��C�*����Z�8[��v�3nV�B,���&�Ϥ^�s���ik��*�H��ў���L���+��|#�e`��k$}�}�Ӭ��ìŶ�$J�?r�}iɅ�*��5���������3���_ƈN�\J�]�f�ef�V�P˭��G��`nE�~%DmQ��P8r����ݿO�����$=Z�o�N�MҢ�Q��s�
��^��V��3�_��~NIs�1*�zj>��jى7�W7!�ui�ݘm(�|2����� B�i�[��s��m=����t:F�߫B��⛤��c��L��T3T�ϫ����R�v)m���?���� Ga��f��H׾��ʭ�)��rk�)J�^o�f��:�F�n�	�H���Ӗ�����ػ�Z6�,la_b�D!��ɑ�5Ы��4o��jHGL�*O�0�����S]������>�~��J��+��"��w�Bg���WS-R�Q�0;gY
�P�O�ܻ�Iyz�ZD�z�aQ�����2k֮(��H�=$������Y��p��@�*���/�ػ�v����"{ƾlj�P0������x0iD� ��e*JW�� ���*eZ������ �v��74�ʟ�Q����N��F��g��p���9�<�ߤ��a�ؙ��Q�!���d������C��CC�$ۼ<cb��V%w��y��yK����u��)�Fuǅ ��O�N�n鿅�r��J$��y�Rՙ/���w$]�	���T�%���Q�߂3�+��s����Sz7]���0ePJ��7ir�0a^�Z�{�!�tE`N�5�+���z�@}�I
����5Ǐ�RW�������V7M�����=�Nh-�dİ�_�(N�Z�E}%|L;�
�h��g
�u�GDV��y@�P�v"�7O��9�~0Q�J���N�h�ӴM�B�8��ۖKU2l�~�n?����\xդ"@h
ކ+D����Xh����[.�=��W�7���r��|#��ja
���6������Y=,��4���;i�?�<�w�\��"Mr�s9�Si,"���v��{�M��Il�\o�S�!�N@z��� �V#���/����qj�d�B7�=n�+���극@7t���������;9	���$���(���M���a%�ۨ��Fs�5}���b��4p@8�5 �����귫І���_b�ث}Pm1���]	�0)︪H��׆��?i�D#�Ǘ�
Q��Y0h<�y��Y�)�SQ^` �����-�Gz��pʺ~�$��6Sw�l���1$ +��zE�eN��b�5��mjA3��f[BL�Kw�F7�*jU ����[ډ0U�-�"0�n�B'�ƣf���=�N	́�Y����D�I1�������:������nN��IZl��N
�?�>��Td)� ��/�*;�"��ͫciA��SlՀ����ی��U�*����*MdM�h�� ����7jh��]S���=�ws��+,�3���/�H�N���&��p��p���ti���
��¿|8���f���@�0���>N�
��O��JC�����8�G#fT~��*�	�C�4?�� m�A;�[�)�_F0n�h�!AT�m^��` �t���r'c��I-��2���?~W�jOi��l+ G���J�ݙ�la�m����p�Aİ��j14{�����,͒`�5�~n"���_��i�����1�,J
��6kp��k�_a|O��S7(�N��h�	��BW�������3�z�L;���q�hq1��)�Т��@ZQ�����Y��0��W��ldG�D�A|��5G�]F6Z�?�f�o��t��2c��>U5��>����_��9�-���%)i+�X�OG�O�Z�P��D'��T"��g�����TxM�b8���٨�*��F�<y�hl�.�-�#�9�J����w���_E|III�}�ity���2��T"rJJe---�����/>8��dvS��"-�(�1�iVI����k54��uQ���)Z�s�5���
�;����l��O�����B�0�.�
�z"�0<�Dl�p������y��F�]�wп�����x�Ȓ�4��d��5��q����P��8���`���0�b\Rol���=?+a���X҅ �u(�F?���8�����_
��bV��j���C�9�]E��{j�8�r�q8���GԴ�������W��;���2f:����;��h��ќ����;UQ��<^�����y���4V��#w�!ײ��2��8�,�����G�T۸;)[���	��ꨈ��ƶG�?*"B�2����֢'�Ջ��v�a����Ш3�Z��|�*��������x���S�V���&Ԋɢ�K�����+��F�bX
1�cc:~P�Ѥ�o_�l�v�&d_����^��^��E��PWJ���+�C��Ȑ�!���1����ii����)��B����Y��ֶ����_d0��B�F�0)֘�J�_�5�9�)�
������`p��7�t.��{{U.\ �p�f����H��U�(��G�����*��D)]Y�sz�B��6��[�w~>��ŋ��W�����yP�1��P����+��i�9�Jî���n�8��{.4E��P�ɷ-��>x\`o��j��~��=�N�� B>&8��"@�J~���_�=�I�2-_nn���V�R��Q�`|�x3�eg{�o�"g`p�3��,O�cU�qS��a&�(��P�D^����^��~�ҫ3�L�0���ٙjM�����R��^�I�|��blwW^���������/�x+�\>�z[̵��!��i;���C��Z�B�$��ح>'ҕ2�Mb�k�c�ga��ԙO���5����+X��D�m��}�h��`�Ì�f�M8[a[娠8/
��)�@���q��&��L(��q��(����maj�/=g��V�����Ԣ�s��^���Ȍ��S����_#"Z��#�AĮ� ������?�~}-+h�ͬ��{Tm��,�8[-$$�z��o����в�c�A��!׸}�5fuC�T���O����m��33<��LN�N�s��=��1�� ��#�������p�Y�߳��1�@u��?�d�N���ER�d�睡��s����E�]ǽ7;��ݼ"�/84�����Ν���Ȁ��L.�ɋ�Q��n14Q�v􉍻���ލ+�i�����FY�y�7������w�{�'��ee�g"Us�֚�����[��B�Y_��K���-�p}��]���JIg]��%<��o̊R;gM���4�^*]��s��i���]����W7�p������h�a��j��=s	Q�шg��ޫ�9T�,��b���8}�[T/��$i|T���VIi	��k|w���Z#�M�&Y*���boo$6J:���;7??2""��˩fܑ?I�a:F!;����ffV�+�L��J`}v���]~���!T��]9�T�	ɢRfFƋ���222&\��Ŵe66>�׫�l�lni�`+G�^��f��i�fuS��cbf��eP�(���������ˡq���9�ȱ�Rq˗�H1��o>�����;+��(�x��"�˃[�𸘘�����TTQ����9�rv�k����=7~1nw��2-�t�f�Д����V9����{e�{ص����h�U�2���bhi�i�X�SpgmQ�m�^AᶒV�%+����ohߡ�@��h���z-�3����O�4%'|�'�{c	�$�!��%��-��.��jVP2]y�o���z���@|Lɻ��X�{ff&q3�*�'�J��X���)�U،"�R�Z����������!��T���d�9r� ���7�����(�H�(UQ���g����v]�qq9�B�����eB�-��y���Ř�_r�/�<9�Ⱦf���z�5�����l����/ �ٳ`��@N�q�q���y�{{.y��9 ߽,����Y�V&�_!:�C���x���t%�Ɔ�L�O��fr��ӭQ;�=�noo��`_�{�����$~�+��"(��5�����W�%�����kS�D����۸a�U@E7�����Ł�+;8S{-{t�Q�Q��ji�|)����P4>�i�?��#�z\� ���d���gfeU��K���,��Cxt���~�vj��IQ�kjh�KAЛ���a�gw�b�V��A�
X0��
S�A�sǰz˃ѡcZ��c
�wl*
�E,rd?T�M�Ё()y���1Y�'W��o�f�T��9�����働t^bb�
/�����
����ڕ��^-� R�4����"$��v,@������x���Y�������Ƈ���Kf��K訠?�`�qe2a(����uQ��4-���W��~��������Cu�o�4*6����,���"��J����-<��Ty�p�r�+墬������BL�/W�*�K1
���=�<�?2�#ޫ�l+Y��t���>{D�/6��%ך
��zV�(?�t��#e�!�B�u�L�5h!�3$�l[�{h]� sM�$el#w��m������4Z���Z����T�0} Y�.��qk������ }��	~P�L1�<AI�uwafc����J?8�P!�=tH�Z'��MC���TUY��>�J����\�2Īƨ��D�	h�_�E~H�
z��ݯ_��dq7T�Օg�>�^@B�룅����?P�ػ�� �����K�?��&��0pY��a@u���,����{�/��Z/�B��>L�mֵ��v�]�.����984����V�B4#�m6�i*�ÔO�p���%�����(Z��$%巶���E��v\������%};I������Dj&}^ ෶X'��+W���vě�<��(����S���L��~��{��1�ˮ�e��W<����dA�*��vrDC�
7|~�� �%�ٽg�_��޷wM�?���/]}u\T]-"�tw�4�H
�)CI*�]"JI�P"%  ��"�tww��w��}����7p�9{?�zֳ�>w��z�u�?g�h�mk~���d�H"Gr�T�?S�YPk�uZ���&����X#Z�av�ve���"����Xw��d�^�:�uu�t��k>̄��
�U��%g�����v_
����]p !f��ى����2��_�?���\��|x.�S�(4=]�C���=���>�%<�
�U(��G?:݁)m*7������vz����|��Eod����2�iXe�#��Zq{ϸ*ٽHHmS�J���N-p�����ЌmM��w:�<��xRE<�|N��j�/�%������U`��*��C(mPߑ_�=���nҶ�����Z�_�!ۄ�/}�"�S	D1	���0��-�B�l�}�at��;�5�J���T�2����QfK�w�C�r��?��}p��g�%�:n��o���h>}���ͽ�X2�Ϛ�j--Mz���f���7�~���r��=��I�583	�Δy�Ejzmgn��Ћ,����|<���Ζp܁��Щ������R�|O��n�f��&�N��n΄k�l�aj�'6h��A��4>"�J�%"#���S�A,r�7��/鴺-y\�''�w�oT��~��E���޾ɼ<�_�?W���!*����/O��%C97y��7|���K����k�~L�҅(e�8m��i���M����r��-�[Ai�$6��k�?]W+M��L���8�/�så=��n}����,u����|��W����E����p�W�i��??Q�/�T6#(��h�ْ�R�JG�;-�����5\�e��ؚHJ���}�7�>V8��!)NlDa�9���3C:�ή�>�/�� � r�@���$�&l�G�ՙTooo�p�ZoW�:C�m��i{�HL�k iw��^b�1o�c�Z
�?��x���92��=U���x����c���P�l�V�tdA��ȝ�$��r�{Mjx����6IQ9�WuurR��~��>������}�S
��`t���!�Hp���A���X��6a���d��H�7�Y�
���$b��y+�����j��D���)��+YLo�Y)!��g����D2w����Q�BF[����/V������t���VO�f��#"���}����8A�T��g�U����#.m�郱�>��@���57��j���Wlͭ�.�6��k�j��ք���o�b�P�Dغi��_�����뀋��J�`�
��*4�N��ъ�:`;o.3R��{�6�Fe���lw�Σ=)�H��1q�yW,���
[�X蠺�+����N���xW�b*��y���h��z�pi����ﺝ�AI�ǳͳԴB'����Mn���n��fx�2U��F�d��I_���Zhq�����*:�#Q4���.パ1�ݭѐ�LQ��)ܜJ���]_�5T��@ 4e�ld	�{���@�?�}I�ؘ��G8ˀ��R������_�� ©���f����h�4�ݓm�����rt���>F�)g�^ (A�BSx �Z��1'��?���ĲM�f��<��VDP�����9��G���?�%)k��r�{�g�(�x�ZS�pKĂ��sC���_�X`�C���ۜ_8��P{���mx�Z&�"�{_�O��5TM����\�`�
�8z^�W��x�0�����l+vrr������b<5�It۪������.��;�}��Z��v�o�\�e���Y[�~+��AXDt~|��fBt�8P�D�6ik�8��<�v�K Vq��T�^�9�z�V��|L��{���d�g�'̿�KtYQ�l��J*�a���ޮ� a��8E�^�B��3 @�� �	�����;L���G��c������gi(���MX�������AT�56�F?qX�z���A��<��%`�3B-y�ż�Q������j��:L���擇:��9�~��z�}�h�ZU���eL=U�{���.��Ff�f��gv���9�6��e:���foD\����CB��f|�N���*���=(O�!�~�>e�c��xQgsp�-Qٓ+,��ǳ|(&�OQR�O��G�ύ���r�q���9)))�' �ń������Y�=��'�:�APf�MBm�P:f���dS*>���6��嶯#��{&��l�L��D�啕� %�+���>�m�:��� ����Ὁ�Y���2s��������VM��Bv�;��Х��"%eeK�7��BAGB�5�	�f..�����L�Ԓ�Nu��u�^�4��gW�������������P̜޲!��Tz�}�ob��+��u�,��9�����:�}dF���g0aL�i��%֬X�ٟ�o�<Bղ��
�����I@F�y^fK�H�, )�V��Pqھ��a�V����-q�Q3�W�m��r)��%=�����#7\K +��94-� !�Jfhm��V4K�����4����'<��C:�m
���B4�J��X]��IJ��/U牚;�kc�d �̒r��X���Ub��̍�i�e�����*�'������F7L��&!��+.�p�yi�= ;$uSY�y�G�*=;j�b���$����2�(�́(�ql�)�����z����L@ 1�ݛ���)G_�����`��~2,�~�S��r��������mB�e�fl�|���Y��MW������fNŌ�2����V��sC��Ĝ��~\1bI�y���C��\��)�"Z%b�F��;oWc�g��#���t*�,�͕D:�H����G�yĮD��W�A�`&ϨO�z��#S�#�������\����W�� �lw����us�_�g����H��i23���9�П���!F�V޿�^��Ʈ����{/�Im��{ҹ�Cs��a�Gv��mZl�7�c5��3Ep�ZdogA��m!����ek�#*B��6|V����Nc��;�ĝ:A�+Zs�Y��p�Ą��	�<`��bdddM[e����m�>��94��T�U�z1��������_�G��x>{~Hʥ��WJ}�;`@iy����~���Ӣ�d����w~����o��X���,p�X���z�IAX���p�痣�?|/ҁq���d��������(��TL�[Ș�`i�6��u��ׇ�V���pݸR�4,��&���a�H!n��ͧp;
�>��2�*��׌

�4�Y�fJ֜�C#_v��Ơ��T�� Q!щm���î�m�*�U��J�-Xs+X��W��ٔ�=�T�4d�Gވ�k�P�Dޒ����(�Gv�=$*Q��tnr?��y�L���dɭ��v��]���k��s��x���׌��l��\C�^�	B��!��d`KPP�N� tXNe�[��M��������}�S�>�|1R�dlt4��w�ߗ�I�ϩp~*{o���Q:�<}|ȳn ��g!c�U}3ө¦&����P;f�ϳ�Hv��6�����A�`�2�3s����^FO�l��}E �6L�~傇������K�~�Sz���1M9$���8� y4��k��Bww���o���ȉ���?�U �[��t��G���e]�2#p�x����S�m<!�	��� �4��'tE�����kmV��;��Q�u`ya3ܝǵY����^�ٱg�lOT��/h/|�<�%��%x1�EQ��N�"a���YU�k͟lt���<��y�`+�c�ː��T�k�����|���USe������	]z�$>4�hfI���"	�W;�"�_����	��Q�j�cD5��������CQ����:b[�r6��r��M�1pw�!���l�a�����[����<�i�� ?V���������[(b8��f]�^�w-���&���Z����3|u��]�WT�����ʈf"%�W9�.t�\i��Ũ��y����oN֗��n�~X_���|ck�������h	�KZ�ռ�n��166P���r�+e9HZ�������:���ubf��?}�MO��3�z#��ж�	%����������
Њ�����e��?��5�O���6��|����#��Xr��EMC���W�7P��5���{"BCS����?)qʮ�$����Z\��@M�@-�����{vE3��gf�gϚ��/��pj*m��\o��K��e�D��i�'�����v��_(;�Ó�׏� ���-T��wQ������>  ]��8���2��nK���Z#Q }�(r��%��rJ��)��|�V�}��	��ѥ��ez;�mS����ώ��w{_�)�7n"����2���j5�sIh��ɯ�|�P�ܕvv�+Y��	���^�����a��Ә�ز<���g�x��SP���́�w4���c��sIa�ج�� -~��*�c�G�Â�Bo����{\&l�ؖ�੝�������V�����]͈�����'n��D��	�ͱ_�""��`���D,�1yr���*>Ni��l�Bڎ�D!�T��05��5�k5/,�Q,����6��D�S@����Q�K\n�p7wq�?dkFpD��ar��4Bd.�P	u������HL��<�T_߀�y&�͑4.�˟�-���ߙ<7ܖL`�滢���Ox��J?xV�HH ;п)è`��{���w��4�+Ft�4(D]����V�wVj��*  ����Ն�'��a-��yԛ�[�#a;;;��� mW	/'��:�� �Ŝk�j(�����d1=:�d�ܷ�[�03$�f�j&��C���3���8^�ޞ�8��ެ���`v\�UM���卽ۓ���pD�~l��g�su瀞4P_W��::fJ(-'�E�F�A�]�/�)����=�������ӝ)<�77�5���iH"u�?�4/8�SΝcd^��� ��uA�q�|s<պ�-��j]dx��ٳ��Uk|���5��d��mҰ�����>0�
�P(l���eb��٬�2���`>a�Ƃ�6qp��R�|T�VHt9���?\gMg���g@�kS�}��|p�G*N.uX�I�H�����Bwq���Kt�a��s^*��*�2
q�Iq)��j���N�$�켼�u�����j��ݽ���=�e����?�~�\b����iļ_%Y���{�y����=A�@dd�s������޴cM�c�h/��H}}}�ggc�������]�����r}����?ha�ꝡq���] ^��a��ެ������5P�ΰC�`�'�@U	t��X�7D��D�Z���~��.fNT"<ѓ�!�@�s���UW}��[9g)�uǺ�r22�����C��C=�zEv��ʽѥN�f���2j��L�� ��o}��g&wu��ֲ�Jo�d�=<�<	e�|)v��ZD�yD{�9"m�
#+��\�r�ϸ�w�
Et����1S6ZT���ڣ����͓�4��DG�R�z*�	D�m�=S�p�%�L3�~��Z�9���)n�< �*�[�T�)�[!����l�ht�>�H����rd�y�&���>A�ޒ�X$@�@%w�zAK�%�h�a���������s4�ڜnh}y	i���/����G��^�]��X��/����2�KV}��8-���Y�RlkYsӪ;2��<����L���Mq�ڿ?������|��t=yX�ˣ�L�7��]&۬�5�Y��5Ȗ����ܸc�ͤ�.����2%$�P�Vi�)f!m�ޚ��~M3�{�1-��ά5�#�]r^#��������D��`�J�X�y�N���A���آVc���qR��8
��c:�Z�P��i������H�9P���>�w�U�Z��_~�}�ts��\DWRj��n�����^2�2���*����4g;��GUp�zw�ߙ1m��}=��ĸx \z=Ǣ������c{ȟާJ�׆���E�*��@C�	����$P/��Bk٤��nkL�4�x��z��q��_������GP< DJ���i#n�i�
����k9���襳?�6�y �"��ōԦ����YN�h%��#�������0�^�_BS�\k�m�6im�("CaҠaa+�,"��	�2�T�,�BS�0�kg�c�
W\$蓙0-��?���;Wnޛ�9}�i��3�'r��uQw����"�\��d4���(�t�D�X݀� ���$9Z,@��&a�0��Hqcr�wE��1@����\�����%j�%b�S���`��%S$-�
���nc��F�}�ހ�ڢ�7h�H'���TY 0�I��N��0ǩ�yq���Ah^��R�5��*�^�:W�IN4,T���!1��}��Lz������E
��
C�R�L��@a������3�³��Z���b[�sO �(i����Bomd���C����9�9e��C��8�k!�W�]̶���K����H����)���ې��BxcU��l���Z\E����
���Mx
s��<b�(�'Q���:�O�c�S�_vH�3;�Q�jA.م�czc>�ﺳx�G�S��V�eAM;eSkQճ���N�"�0U��6ʬ����t�RGE���n�@���8���d�k�eZ"3�����ŝ�{Pf�z#7*��T]�Rf5���
�N�Yd�TzuX��
V�y8�F�.��w�dК��{dkHttt�����j���݀�b�'XX�s1�d�����0��54�It���TהԪ�	��f���g���S�R�ܣ�,�i��+i\����I���ճt�EPÅ?u'���*���ʖ����u�v��ߺL�i�Ԅ�O��ќr��gN�ecv�*�
n$���xR�Y�dr�>�_�"���d�\WMT�J,���i��|��K�·h�Y�c�w��z�	-�z��wM����ch� �k=�g��~"/V$�=��/N;P�E��|�R��tG,�N�@U�X��u{#_��E%�5:sQ���6+].��cU�
vA� �a7>fm���n��~�B����]ה.�!�y��w��w"fMC@��Z|��M�1��޲)�T�����H�1���Oi�g����r*�6��'�O�M�Jw]&�~,��˿h�zΥ�mE�Cz"�B$��������Mn�"��?Mi�â=c�J�fҬ_�n*�p���� `|�jNX��Gv{�摙$q-w����h�[����f��2\L�q�]!%��r1�:�U%� 밧����ˤ(͜P�������w
��s�dz��zf���O�����4VKq3�b-V�N��hߣ,�B�UH,��6i�>`��ט�sL�z!V�RgW���m,M,c
U2|-E�����	�1U�$!U�sŗ�tr�KwK�+�6�Ϸ���ې�cdF'�G��O[$MwiOȫ̬ʴLC�ph���t{"W�""BAy?��^����E/샳%�B�6��=<�	N�=O-�CtJcȉI�+P�n{�{�V��^SI��.��֍3��m�U+"���,5�	N�98o;ɯ,������#��U]��k�h:�2�Vr���^�uO����*�T�R��ˏ_��M� ����\Dzo��E�U�p7jѢ�D�Y�B�g����^��D�J��fO�u����]{"�a�ܴB�~H���MH��jI��뤣آN��4Us�b�f��`��9?4������W��m��4ʇz"�2�����bi�
U5t�9>_��*�b�&h�W��nzR.�:�4D���?F�!�ԛ�V��yo��ĵ/1��$}B����<o�}|�m��:�
�t�Ħ�mJ���b*��O�|��Ut,n�#�?Y���	�L�ɯG&�9�YM~��6�cv�@�B�����z���� ��f�c{��m��Ͷ��170�j�}�OD��O��o\�MplmS�.�勬�o���P6��'{yox�{������(��Z�.�u�z�s?Qd��TW[�N�������p�Bp�q�W��Tv�H/�m�����D22�9ѵ����&Q�X�mBoFs�X��*J ��^I�23ۀ���P��8�z%&��@�\�o���]�_� x�&��G���i�����J6*�w!���1���ә>R�޼mbK��:m�]>�Ҍ^4��:_#	��tC.�����P�db%�*��5���ǥ�`%��B�7�����c�ۯ�̭_?Q�]ŗR� ]���xP����B�߫z"�ˬ"mL����~T�MwII\����9�n^���?F��� ��ݙ�o1�VN�V�6>�B��m��������&�3'5��k�i�왕���4)vmH�
3)���Z�5�g�F�2���+)�+�Ӊ|�3�o8e�Z-�3p���s6J�#&�z�ٖ�B>f�֏�u��gI>fI�SS� ��u&�(�N���s��M��|{�	��HW��_����a�<��0�>w)F)�g��B5�xw|�&�������M�rV:�~O�iv̜�N�;��I	�(E��bTp��p_=��z�iJ���]lؑ��޳�V7�k�����{��#��� '�mJ���F��`�`1؃ׇ7ח���R:��;v�Z�Ab4k�=��6�3�w�~"�L���/�y�f67���ÂB�+&9���{S9�B��{]+3bq��1B�xC�ߏ�cx�˺�ٺ���X
t�
�ܺ��uJJ��L���QyQ�mr.W�*\9��}2��(2�n�w��ݙ
��vcG�_7ڑʿ���D��̢X�U�+I�����_��S�|9�Nd�3J���
~����Z����� a*�$����[(�����$],�~:ř��~|rِ@��O�%Il%�����C�EJ&��B���NBx�)�VS]�DKi~��c(m~�� �Ĉ�9q+'b�$'��ن�-`�	�����d����yS�ǚ�S@�ʽ��c=}S,PB(�5&�^]��1v�_u&���dd�I�i���Ӻ·$!�d�.�q�.�j.���,ۨ�d�U��C�Q��?�q3�Zo`r�0��/�����|��)M��t\��B�c$�.Q.ͦ�d�6i�z|r��<��-څ�-j�~�fe�VUxs�S{B]c�����������\�G��#�1���3�����H#���7F+�=�Lʲ�jl��/�572��\�.7�N������!�ZD[[�?Jw%�'_�!��)0)���>Sb�䎒bJ�����)O&�I�
��c�WrG���,�i^Jh1C�I(�bQ7!�|�F��Z�*h��5��n�����}���w
6K�����s��i�@�'�߽�_�\����'�DQ��D�K�I�JD�xI�<�~4�F��=�7O֑��l{�B�PO;;vdD�,���5�%(v�HapL�M�8�Z��\�}������!����xy<M�R������a�������"*
	X�оNLN~B{��x%��Ww��7pt��(���8
��(`���	��y!7����{�O�~��ǋD��K���멽���$Sin���]��Ck͇�cJ�6� L���rA��c,т}Q�9;�����2�\��t�+���?1��e7/'�����fTr�1����tJ����iE���8�{f���v�]1���c�5��9�)��"\��GıL�'�m������]�M��d�w���{�nO�I�p���d>�������:r�f��1���քK�Nn�ԉ�)�UCib�����,�/��1�Bsw\뉬��%�$AX�V!���cʗa��| �Q�ѯ�!��/)���W|�����L��� ]��w�uO��yWz#�Ƚ����v��VF̊�N��� Z����G�y�X ����g�lX�&O�HR�:p:�ݻ@���O�R�e>rj��)��?���G������*��"��h7�>���R􊨷��/�~��d�UЯ��D��B�Vx�@�G�ٝ��
�@.��]���Lv�Dl��{,,�%������G�!�B�~+I�`���S�wg���uvٸ*������ڃ��9m�he�wL����O'�N��HT�A��8��죞�{�!t�������!k4n9?���,���Z3�À�_�}Ԝ��U��o�?�H�!��$���x��-m��A?�"�ݟ�+ʪɔJ���PK   �}Xa6�~  y     jsons/user_defined.json��]O�8��
�u��N�vv��Ѱp�B#�q ���|B���NR����a�u��8�y}Λ��{ܚh��i�g&/*�E��iڢ���ّ�O�[�h���˟3u7�]5Y_T���ٹ�Q����ͣ�1:-tS�ꚺ,M]/�@�]�e���,����0�RF!�1�(�S SbG���ulL��b�M�|�Zh�?�8��e�h� ��H�	 ��FS̴񶺱���t ����G���^��q����)���M�nK����vXk3{�����aG��i�����튪��k
�n�pC���O�Ҏ ����BѮ*}[7vJ���nM�R3�uyvy�e=/����y�n�_���߾���b˂��Lk:/��X�%1��R�KAT�g2�)����_w����
�a�ʎ��҅� �
z����(�=��ߕ���C]Q��_?ԕ���C]A��_1?��S���B/�'~ꌢ` v��cg4�°�C re�p��X�+,D°t �\m!���-����-���/x�h�@l���,H�~������
?��F�T�A�����E���.H��ϔ.H�����.H����/H�ں�ؿ'o�P4�Y��l+?5ؚN%�@KF%2)�����+�3B�]��m�i�bgv~��j{��C�m��v���]%�C��g�v�m�p^����^�h��4?�sߏ��a{|U��Jw}c��^�����v��RW��^���x�n�Im}�d^J������5��|k�N֛�c�>��w��.���N]������Nsh�1H)�@r�3�#���f�ƞM$�q1�,�`�R`�*����aIY� ������E�HN��6�ΤF) �$ �	L0ɍH�ˤ���WC1BH�9��D�%L�'\��0�:���Ĉ�<l�6�	�_����E���`3r/
�04���ϛ��ڕ�׿�NM7�y_#�ն�Oӻ�"��0�@e�"�� ����4�*�� ��B:J	(K)P9I ��J��P�lw0~>�%�Y��&�MiS��'>DHd�J&9Z0�cf���G���R�/$�^n�G���o��� IX�Q�!	�ra&	D���5'(��i.��:���{��1K����PK
   �}XG��   �Y                   cirkitFile.jsonPK
   JrX �/��  �  /             M  images/25830125-c098-459c-a621-2bf82c8cd0ac.pngPK
   }X�_B�   #  /             .  images/530fdb4e-21ab-4901-ad86-29119845d103.jpgPK
   }Xv��^}%  �)  /             Y4  images/b7b52948-3c4e-4eaa-8c83-bc90923fe796.jpgPK
   �}X$7h�!  �!  /             #Z  images/c6364832-c854-438f-b38b-75bf2a0cd33f.pngPK
   JrXPD> �  ��  /             f|  images/ee20a1cf-a7e8-45b4-af39-6cac45e8073d.pngPK
   �}XP��/�  ǽ  /             �\ images/f42d805d-3c79-4d19-85d7-77e6ec425ca7.pngPK
   �}Xa6�~  y               % jsons/user_defined.jsonPK      �  �   